`ifndef MAIN_RFG_PKG
`define MAIN_RFG_PKG
package main_rfg_pkg;
    enum {
    SCRATCHPAD0 = 8'h0,
    SCRATCHPAD1 = 8'h1
    } addresses;
endpackage
`endif
