VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO COMP_R2RV2_BIAS
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN COMP_R2RV2_BIAS 0 0 ;
  SIZE 37.66 BY 30.18 ;
  SYMMETRY X Y R90 ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER ME4 ;
        RECT 2.9 25.87 34.76 28.18 ;
        RECT 32.76 2 34.76 28.18 ;
        RECT 2.9 2 34.76 4.31 ;
        RECT 22.72 25.06 23.37 28.18 ;
        RECT 7.41 25.1 7.79 28.18 ;
        RECT 2.9 9.83 5.67 10.81 ;
        RECT 2.9 2 4.9 28.18 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER ME3 ;
        RECT 0.9 28.18 36.76 30.18 ;
        RECT 34.76 0 36.76 30.18 ;
        RECT 31.1 24.06 36.76 24.44 ;
        RECT 0.9 0 36.76 2 ;
        RECT 31.42 0 31.92 5.33 ;
        RECT 0.9 5.13 7.29 5.63 ;
        RECT 0.9 19.12 5.58 20.12 ;
        RECT 0.9 0 2.9 30.18 ;
    END
  END VDD
  PIN VREF
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 0 12.8 0.59 13.39 ;
    END
  END VREF
  PIN VOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 37.16 14.22 37.66 14.72 ;
    END
  END VOUT
  PIN VIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 0 13.89 0.55 14.44 ;
    END
  END VIN2
  PIN VIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 0 14.74 0.55 15.29 ;
    END
  END VIN1
  OBS
    LAYER ME1 ;
      RECT 30.83 14.22 37.66 14.72 ;
    LAYER ME1 SPACING 0.09 ;
      RECT 1 1 36.66 29.18 ;
      RECT 1 14.22 37.66 14.72 ;
      RECT 0 12.86 0.5 13.36 ;
      RECT 0 13.91 0.5 14.41 ;
      RECT 0 14.76 0.5 15.26 ;
    LAYER VI1 SPACING 0.1 ;
      RECT 37.48 14.32 37.58 14.42 ;
      RECT 37.48 14.52 37.58 14.62 ;
      RECT 37.24 14.32 37.34 14.42 ;
      RECT 37.24 14.52 37.34 14.62 ;
      RECT 1 1 36.66 29.18 ;
      RECT 0.32 12.96 0.42 13.06 ;
      RECT 0.32 13.16 0.42 13.26 ;
      RECT 0.32 14.01 0.42 14.11 ;
      RECT 0.32 14.21 0.42 14.31 ;
      RECT 0.32 14.86 0.42 14.96 ;
      RECT 0.32 15.06 0.42 15.16 ;
      RECT 0.08 12.96 0.18 13.06 ;
      RECT 0.08 13.16 0.18 13.26 ;
      RECT 0.08 14.01 0.18 14.11 ;
      RECT 0.08 14.21 0.18 14.31 ;
      RECT 0.08 14.86 0.18 14.96 ;
      RECT 0.08 15.06 0.18 15.16 ;
    LAYER ME2 ;
      RECT 0.85 13.89 5.79 14.44 ;
      RECT 0.85 14.74 5.79 15.29 ;
      RECT 0.89 12.8 0.9 13.39 ;
    LAYER ME2 SPACING 0.1 ;
      RECT 1 1 36.66 29.18 ;
      RECT 0.73 14.74 36.66 15.29 ;
      RECT 0.73 13.89 36.66 14.44 ;
      RECT 0.77 12.8 0.9 13.39 ;
    LAYER VI2 SPACING 0.1 ;
      RECT 37.48 14.32 37.58 14.42 ;
      RECT 37.48 14.52 37.58 14.62 ;
      RECT 37.24 14.32 37.34 14.42 ;
      RECT 37.24 14.52 37.34 14.62 ;
      RECT 1 1 36.66 29.18 ;
      RECT 0.32 12.96 0.42 13.06 ;
      RECT 0.32 13.16 0.42 13.26 ;
      RECT 0.32 14.01 0.42 14.11 ;
      RECT 0.32 14.21 0.42 14.31 ;
      RECT 0.32 14.86 0.42 14.96 ;
      RECT 0.32 15.06 0.42 15.16 ;
      RECT 0.08 12.96 0.18 13.06 ;
      RECT 0.08 13.16 0.18 13.26 ;
      RECT 0.08 14.01 0.18 14.11 ;
      RECT 0.08 14.21 0.18 14.31 ;
      RECT 0.08 14.86 0.18 14.96 ;
      RECT 0.08 15.06 0.18 15.16 ;
    LAYER ME3 SPACING 0.1 ;
      RECT 3.08 24.62 34.58 28 ;
      RECT 3.08 20.3 30.92 28 ;
      RECT 32.1 2.18 34.58 23.88 ;
      RECT 5.76 5.81 34.58 23.88 ;
      RECT 7.47 5.51 34.58 23.88 ;
      RECT 3.08 5.81 34.58 18.94 ;
      RECT 7.47 2.18 31.24 23.88 ;
      RECT 3.08 2.18 31.24 4.95 ;
      RECT 37.16 14.22 37.66 14.72 ;
      RECT 0 12.86 0.5 13.36 ;
      RECT 0 13.91 0.5 14.41 ;
      RECT 0 14.76 0.5 15.26 ;
    LAYER VI3 SPACING 0.1 ;
      RECT 37.48 14.32 37.58 14.42 ;
      RECT 37.48 14.52 37.58 14.62 ;
      RECT 37.24 14.32 37.34 14.42 ;
      RECT 37.24 14.52 37.34 14.62 ;
      RECT 1 1 36.66 29.18 ;
      RECT 0.32 12.96 0.42 13.06 ;
      RECT 0.32 13.16 0.42 13.26 ;
      RECT 0.32 14.01 0.42 14.11 ;
      RECT 0.32 14.21 0.42 14.31 ;
      RECT 0.32 14.86 0.42 14.96 ;
      RECT 0.32 15.06 0.42 15.16 ;
      RECT 0.08 12.96 0.18 13.06 ;
      RECT 0.08 13.16 0.18 13.26 ;
      RECT 0.08 14.01 0.18 14.11 ;
      RECT 0.08 14.21 0.18 14.31 ;
      RECT 0.08 14.86 0.18 14.96 ;
      RECT 0.08 15.06 0.18 15.16 ;
    LAYER ME4 SPACING 0.1 ;
      RECT 23.55 24.62 32.58 25.69 ;
      RECT 7.97 4.49 22.54 25.69 ;
      RECT 5.08 20.3 7.23 25.69 ;
      RECT 5.08 20.3 22.54 24.92 ;
      RECT 7.47 4.49 30.92 24.88 ;
      RECT 32.1 4.49 32.58 23.88 ;
      RECT 5.76 10.99 32.58 23.88 ;
      RECT 7.47 5.51 32.58 23.88 ;
      RECT 5.08 10.99 32.58 18.94 ;
      RECT 5.85 5.81 32.58 23.88 ;
      RECT 5.08 5.81 32.58 9.65 ;
      RECT 7.47 4.49 31.24 23.88 ;
      RECT 5.08 4.49 31.24 4.95 ;
      RECT 37.16 14.22 37.66 14.72 ;
      RECT 0 12.86 0.5 13.36 ;
      RECT 0 13.91 0.5 14.41 ;
      RECT 0 14.76 0.5 15.26 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END COMP_R2RV2_BIAS

MACRO DACR2R_8BITV1_PWRRING
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DACR2R_8BITV1_PWRRING 0 0 ;
  SIZE 601.85 BY 183.81 ;
  SYMMETRY X Y R90 ;
  PIN dac[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 48.8 0 49.4 0.6 ;
    END
  END dac[0]
  PIN dac[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 117.6 0 118.2 0.6 ;
    END
  END dac[1]
  PIN dac[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 186.5 0 187.1 0.6 ;
    END
  END dac[2]
  PIN dac[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 255.4 0 256 0.6 ;
    END
  END dac[3]
  PIN dac[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 324.1 0 324.7 0.6 ;
    END
  END dac[4]
  PIN dac[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 393 0 393.6 0.6 ;
    END
  END dac[5]
  PIN dac[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 461.7 0 462.3 0.6 ;
    END
  END dac[6]
  PIN dac[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 530.6 0 531.2 0.6 ;
    END
  END dac[7]
  PIN dacout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 598.66 0 599.16 0.5 ;
    END
  END dacout
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER ME3 ;
        RECT 0 181.81 601.85 183.81 ;
        RECT 599.85 0.9 601.85 183.81 ;
        RECT 0 0.9 601.85 2.9 ;
        RECT 38.6 0.9 39.71 6.9 ;
        RECT 0 0.9 2 183.81 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER ME4 ;
        RECT 2 179.5 599.85 181.81 ;
        RECT 597.85 2.9 599.85 181.81 ;
        RECT 2 2.9 599.85 5.21 ;
        RECT 2 2.9 4 181.81 ;
    END
  END GND
  OBS
    LAYER ME1 SPACING 0.09 ;
      RECT 1 1 600.85 182.81 ;
      RECT 598.66 0 599.16 0.5 ;
      RECT 530.61 0 531.11 0.5 ;
      RECT 461.78 0 462.28 0.5 ;
      RECT 393.05 0 393.55 0.5 ;
      RECT 324.12 0 324.62 0.5 ;
      RECT 255.49 0 255.99 0.5 ;
      RECT 186.56 0 187.06 0.5 ;
      RECT 117.63 0 118.13 0.5 ;
      RECT 48.84 0 49.34 0.5 ;
    LAYER VI1 SPACING 0.1 ;
      RECT 1 1 600.85 182.81 ;
      RECT 598.98 0.1 599.08 0.2 ;
      RECT 598.98 0.3 599.08 0.4 ;
      RECT 598.74 0.1 598.84 0.2 ;
      RECT 598.74 0.3 598.84 0.4 ;
      RECT 530.93 0.1 531.03 0.2 ;
      RECT 530.93 0.3 531.03 0.4 ;
      RECT 530.69 0.1 530.79 0.2 ;
      RECT 530.69 0.3 530.79 0.4 ;
      RECT 462.1 0.1 462.2 0.2 ;
      RECT 462.1 0.3 462.2 0.4 ;
      RECT 461.86 0.1 461.96 0.2 ;
      RECT 461.86 0.3 461.96 0.4 ;
      RECT 393.37 0.1 393.47 0.2 ;
      RECT 393.37 0.3 393.47 0.4 ;
      RECT 393.13 0.1 393.23 0.2 ;
      RECT 393.13 0.3 393.23 0.4 ;
      RECT 324.44 0.1 324.54 0.2 ;
      RECT 324.44 0.3 324.54 0.4 ;
      RECT 324.2 0.1 324.3 0.2 ;
      RECT 324.2 0.3 324.3 0.4 ;
      RECT 255.81 0.1 255.91 0.2 ;
      RECT 255.81 0.3 255.91 0.4 ;
      RECT 255.57 0.1 255.67 0.2 ;
      RECT 255.57 0.3 255.67 0.4 ;
      RECT 186.88 0.1 186.98 0.2 ;
      RECT 186.88 0.3 186.98 0.4 ;
      RECT 186.64 0.1 186.74 0.2 ;
      RECT 186.64 0.3 186.74 0.4 ;
      RECT 117.95 0.1 118.05 0.2 ;
      RECT 117.95 0.3 118.05 0.4 ;
      RECT 117.71 0.1 117.81 0.2 ;
      RECT 117.71 0.3 117.81 0.4 ;
      RECT 49.16 0.1 49.26 0.2 ;
      RECT 49.16 0.3 49.26 0.4 ;
      RECT 48.92 0.1 49.02 0.2 ;
      RECT 48.92 0.3 49.02 0.4 ;
    LAYER ME2 ;
      RECT 598.69 0.8 599.14 11.53 ;
      RECT 530.6 0.9 531.2 5.1 ;
      RECT 461.7 0.9 462.3 5.1 ;
      RECT 393 0.9 393.6 5.1 ;
      RECT 324.1 0.9 324.7 5.1 ;
      RECT 255.4 0.9 256 5.1 ;
      RECT 186.5 0.9 187.1 5.1 ;
      RECT 117.6 0.9 118.2 5.1 ;
      RECT 48.8 0.9 49.4 5.1 ;
    LAYER ME2 SPACING 0.1 ;
      RECT 1 1 600.85 182.81 ;
      RECT 598.69 0.68 599.14 182.81 ;
      RECT 530.6 0.78 531.2 182.81 ;
      RECT 461.7 0.78 462.3 182.81 ;
      RECT 393 0.78 393.6 182.81 ;
      RECT 324.1 0.78 324.7 182.81 ;
      RECT 255.4 0.78 256 182.81 ;
      RECT 186.5 0.78 187.1 182.81 ;
      RECT 117.6 0.78 118.2 182.81 ;
      RECT 48.8 0.78 49.4 182.81 ;
    LAYER VI2 SPACING 0.1 ;
      RECT 1 1 600.85 182.81 ;
      RECT 598.98 0.1 599.08 0.2 ;
      RECT 598.98 0.3 599.08 0.4 ;
      RECT 598.74 0.1 598.84 0.2 ;
      RECT 598.74 0.3 598.84 0.4 ;
      RECT 530.93 0.1 531.03 0.2 ;
      RECT 530.93 0.3 531.03 0.4 ;
      RECT 530.69 0.1 530.79 0.2 ;
      RECT 530.69 0.3 530.79 0.4 ;
      RECT 462.1 0.1 462.2 0.2 ;
      RECT 462.1 0.3 462.2 0.4 ;
      RECT 461.86 0.1 461.96 0.2 ;
      RECT 461.86 0.3 461.96 0.4 ;
      RECT 393.37 0.1 393.47 0.2 ;
      RECT 393.37 0.3 393.47 0.4 ;
      RECT 393.13 0.1 393.23 0.2 ;
      RECT 393.13 0.3 393.23 0.4 ;
      RECT 324.44 0.1 324.54 0.2 ;
      RECT 324.44 0.3 324.54 0.4 ;
      RECT 324.2 0.1 324.3 0.2 ;
      RECT 324.2 0.3 324.3 0.4 ;
      RECT 255.81 0.1 255.91 0.2 ;
      RECT 255.81 0.3 255.91 0.4 ;
      RECT 255.57 0.1 255.67 0.2 ;
      RECT 255.57 0.3 255.67 0.4 ;
      RECT 186.88 0.1 186.98 0.2 ;
      RECT 186.88 0.3 186.98 0.4 ;
      RECT 186.64 0.1 186.74 0.2 ;
      RECT 186.64 0.3 186.74 0.4 ;
      RECT 117.95 0.1 118.05 0.2 ;
      RECT 117.95 0.3 118.05 0.4 ;
      RECT 117.71 0.1 117.81 0.2 ;
      RECT 117.71 0.3 117.81 0.4 ;
      RECT 49.16 0.1 49.26 0.2 ;
      RECT 49.16 0.3 49.26 0.4 ;
      RECT 48.92 0.1 49.02 0.2 ;
      RECT 48.92 0.3 49.02 0.4 ;
    LAYER ME3 SPACING 0.1 ;
      RECT 2.18 7.08 599.67 181.63 ;
      RECT 39.89 3.08 599.67 181.63 ;
      RECT 2.18 3.08 38.42 181.63 ;
      RECT 598.66 0 599.16 0.5 ;
      RECT 530.61 0 531.11 0.5 ;
      RECT 461.78 0 462.28 0.5 ;
      RECT 393.05 0 393.55 0.5 ;
      RECT 324.12 0 324.62 0.5 ;
      RECT 255.49 0 255.99 0.5 ;
      RECT 186.56 0 187.06 0.5 ;
      RECT 117.63 0 118.13 0.5 ;
      RECT 48.84 0 49.34 0.5 ;
    LAYER VI3 SPACING 0.1 ;
      RECT 1 1 600.85 182.81 ;
      RECT 598.98 0.1 599.08 0.2 ;
      RECT 598.98 0.3 599.08 0.4 ;
      RECT 598.74 0.1 598.84 0.2 ;
      RECT 598.74 0.3 598.84 0.4 ;
      RECT 530.93 0.1 531.03 0.2 ;
      RECT 530.93 0.3 531.03 0.4 ;
      RECT 530.69 0.1 530.79 0.2 ;
      RECT 530.69 0.3 530.79 0.4 ;
      RECT 462.1 0.1 462.2 0.2 ;
      RECT 462.1 0.3 462.2 0.4 ;
      RECT 461.86 0.1 461.96 0.2 ;
      RECT 461.86 0.3 461.96 0.4 ;
      RECT 393.37 0.1 393.47 0.2 ;
      RECT 393.37 0.3 393.47 0.4 ;
      RECT 393.13 0.1 393.23 0.2 ;
      RECT 393.13 0.3 393.23 0.4 ;
      RECT 324.44 0.1 324.54 0.2 ;
      RECT 324.44 0.3 324.54 0.4 ;
      RECT 324.2 0.1 324.3 0.2 ;
      RECT 324.2 0.3 324.3 0.4 ;
      RECT 255.81 0.1 255.91 0.2 ;
      RECT 255.81 0.3 255.91 0.4 ;
      RECT 255.57 0.1 255.67 0.2 ;
      RECT 255.57 0.3 255.67 0.4 ;
      RECT 186.88 0.1 186.98 0.2 ;
      RECT 186.88 0.3 186.98 0.4 ;
      RECT 186.64 0.1 186.74 0.2 ;
      RECT 186.64 0.3 186.74 0.4 ;
      RECT 117.95 0.1 118.05 0.2 ;
      RECT 117.95 0.3 118.05 0.4 ;
      RECT 117.71 0.1 117.81 0.2 ;
      RECT 117.71 0.3 117.81 0.4 ;
      RECT 49.16 0.1 49.26 0.2 ;
      RECT 49.16 0.3 49.26 0.4 ;
      RECT 48.92 0.1 49.02 0.2 ;
      RECT 48.92 0.3 49.02 0.4 ;
    LAYER ME4 SPACING 0.1 ;
      RECT 4.18 7.08 597.67 179.32 ;
      RECT 39.89 5.39 597.67 179.32 ;
      RECT 4.18 5.39 38.42 179.32 ;
      RECT 598.66 0 599.16 0.5 ;
      RECT 530.61 0 531.11 0.5 ;
      RECT 461.78 0 462.28 0.5 ;
      RECT 393.05 0 393.55 0.5 ;
      RECT 324.12 0 324.62 0.5 ;
      RECT 255.49 0 255.99 0.5 ;
      RECT 186.56 0 187.06 0.5 ;
      RECT 117.63 0 118.13 0.5 ;
      RECT 48.84 0 49.34 0.5 ;
  END
  PROPERTY CatenaDesignType "chipAssembly" ;
END DACR2R_8BITV1_PWRRING

MACRO OSC_RINGTOPV1_NOVAR
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN OSC_RINGTOPV1_NOVAR 0 0 ;
  SIZE 102 BY 39.9 ;
  SYMMETRY X Y R90 ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER ME4 ;
        RECT 2 35.59 100 37.9 ;
        RECT 98 2.9 100 37.9 ;
        RECT 2 2.9 100 5.21 ;
        RECT 2 2.9 4 37.9 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER ME3 ;
        RECT 0 37.9 102 39.9 ;
        RECT 100 0.65 102 39.9 ;
        RECT 0.01 0.65 102 2.65 ;
        RECT 0 0.9 2 39.9 ;
    END
  END VDD
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME2 ;
        RECT 82.04 0 82.54 0.5 ;
    END
  END EN
  PIN CKOUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER ME1 ;
        RECT 91.66 0 92.16 0.5 ;
    END
  END CKOUT
  OBS
    LAYER ME1 ;
      RECT 91.8 0.8 92.01 9.31 ;
      RECT 80.78 18.94 81.28 39.9 ;
      RECT 62.52 33.65 63.79 39.89 ;
      RECT 58.46 31.98 59.05 39.9 ;
      RECT 0 5.61 4.73 5.88 ;
      RECT 0 10.34 4.73 10.61 ;
    LAYER ME1 SPACING 0.09 ;
      RECT 80.78 1 81.28 39.9 ;
      RECT 58.46 1 59.05 39.9 ;
      RECT 62.52 1 63.79 39.89 ;
      RECT 1 1 101 38.9 ;
      RECT 0 10.34 101 10.61 ;
      RECT 0 5.61 101 5.88 ;
      RECT 91.8 0.67 92.01 38.9 ;
      RECT 82.04 0 82.54 0.5 ;
    LAYER VI1 SPACING 0.1 ;
      RECT 81.1 1 81.2 39.05 ;
      RECT 80.86 1 80.96 39.05 ;
      RECT 58.915 1 59.015 38.95 ;
      RECT 58.705 1 58.805 38.95 ;
      RECT 58.495 1 58.595 38.95 ;
      RECT 63.63 1 63.73 38.945 ;
      RECT 63.42 1 63.52 38.945 ;
      RECT 63.21 1 63.31 38.945 ;
      RECT 63 1 63.1 38.945 ;
      RECT 62.79 1 62.89 38.945 ;
      RECT 62.58 1 62.68 38.945 ;
      RECT 1 1 101 38.9 ;
      RECT 0.85 10.42 101 10.52 ;
      RECT 0.85 5.69 101 5.79 ;
      RECT 91.98 0.1 92.08 0.2 ;
      RECT 91.98 0.3 92.08 0.4 ;
      RECT 91.74 0.1 91.84 0.2 ;
      RECT 91.74 0.3 91.84 0.4 ;
      RECT 82.36 0.1 82.46 0.2 ;
      RECT 82.36 0.3 82.46 0.4 ;
      RECT 82.12 0.1 82.22 0.2 ;
      RECT 82.12 0.3 82.22 0.4 ;
      RECT 81.1 39.15 81.2 39.25 ;
      RECT 81.1 39.35 81.2 39.45 ;
      RECT 81.1 39.55 81.2 39.65 ;
      RECT 81.1 39.75 81.2 39.85 ;
      RECT 80.86 39.15 80.96 39.25 ;
      RECT 80.86 39.35 80.96 39.45 ;
      RECT 80.86 39.55 80.96 39.65 ;
      RECT 80.86 39.75 80.96 39.85 ;
      RECT 63.63 39.055 63.73 39.155 ;
      RECT 63.63 39.265 63.73 39.365 ;
      RECT 63.63 39.475 63.73 39.575 ;
      RECT 63.63 39.685 63.73 39.785 ;
      RECT 63.42 39.055 63.52 39.155 ;
      RECT 63.42 39.265 63.52 39.365 ;
      RECT 63.42 39.475 63.52 39.575 ;
      RECT 63.42 39.685 63.52 39.785 ;
      RECT 63.21 39.055 63.31 39.155 ;
      RECT 63.21 39.265 63.31 39.365 ;
      RECT 63.21 39.475 63.31 39.575 ;
      RECT 63.21 39.685 63.31 39.785 ;
      RECT 63 39.055 63.1 39.155 ;
      RECT 63 39.265 63.1 39.365 ;
      RECT 63 39.475 63.1 39.575 ;
      RECT 63 39.685 63.1 39.785 ;
      RECT 62.79 39.055 62.89 39.155 ;
      RECT 62.79 39.265 62.89 39.365 ;
      RECT 62.79 39.475 62.89 39.575 ;
      RECT 62.79 39.685 62.89 39.785 ;
      RECT 62.58 39.055 62.68 39.155 ;
      RECT 62.58 39.265 62.68 39.365 ;
      RECT 62.58 39.475 62.68 39.575 ;
      RECT 62.58 39.685 62.68 39.785 ;
      RECT 58.915 39.06 59.015 39.16 ;
      RECT 58.915 39.27 59.015 39.37 ;
      RECT 58.915 39.48 59.015 39.58 ;
      RECT 58.915 39.69 59.015 39.79 ;
      RECT 58.705 39.06 58.805 39.16 ;
      RECT 58.705 39.27 58.805 39.37 ;
      RECT 58.705 39.48 58.805 39.58 ;
      RECT 58.705 39.69 58.805 39.79 ;
      RECT 58.495 39.06 58.595 39.16 ;
      RECT 58.495 39.27 58.595 39.37 ;
      RECT 58.495 39.48 58.595 39.58 ;
      RECT 58.495 39.69 58.595 39.79 ;
    LAYER ME2 ;
      RECT 89.37 33.76 90.37 39.9 ;
      RECT 82.2 0.8 82.4 6.92 ;
      RECT 80.78 37.9 81.28 39.9 ;
      RECT 62.52 37.9 63.79 39.89 ;
      RECT 58.46 37.9 59.05 39.9 ;
      RECT 0.82 5.66 1.18 5.82 ;
      RECT 0.82 10.39 1.18 10.55 ;
    LAYER ME2 SPACING 0.1 ;
      RECT 89.37 1 90.37 39.9 ;
      RECT 80.78 1 81.28 39.9 ;
      RECT 58.46 1 59.05 39.9 ;
      RECT 62.52 1 63.79 39.89 ;
      RECT 1 1 101 38.9 ;
      RECT 0.82 10.39 101 10.55 ;
      RECT 0.82 5.66 101 5.82 ;
      RECT 82.2 0.68 82.4 38.9 ;
      RECT 91.66 0 92.16 0.5 ;
    LAYER VI2 SPACING 0.1 ;
      RECT 81.1 1 81.2 39.05 ;
      RECT 80.86 1 80.96 39.05 ;
      RECT 90.24 1 90.34 38.95 ;
      RECT 90.03 1 90.13 38.95 ;
      RECT 89.82 1 89.92 38.95 ;
      RECT 89.61 1 89.71 38.95 ;
      RECT 89.4 1 89.5 38.95 ;
      RECT 58.915 1 59.015 38.95 ;
      RECT 58.705 1 58.805 38.95 ;
      RECT 58.495 1 58.595 38.95 ;
      RECT 63.63 1 63.73 38.945 ;
      RECT 63.42 1 63.52 38.945 ;
      RECT 63.21 1 63.31 38.945 ;
      RECT 63 1 63.1 38.945 ;
      RECT 62.79 1 62.89 38.945 ;
      RECT 62.58 1 62.68 38.945 ;
      RECT 1 1 101 38.9 ;
      RECT 0.85 10.42 101 10.52 ;
      RECT 0.85 5.69 101 5.79 ;
      RECT 91.98 0.1 92.08 0.2 ;
      RECT 91.98 0.3 92.08 0.4 ;
      RECT 91.74 0.1 91.84 0.2 ;
      RECT 91.74 0.3 91.84 0.4 ;
      RECT 90.24 39.06 90.34 39.16 ;
      RECT 90.24 39.27 90.34 39.37 ;
      RECT 90.24 39.48 90.34 39.58 ;
      RECT 90.24 39.69 90.34 39.79 ;
      RECT 90.03 39.06 90.13 39.16 ;
      RECT 90.03 39.27 90.13 39.37 ;
      RECT 90.03 39.48 90.13 39.58 ;
      RECT 90.03 39.69 90.13 39.79 ;
      RECT 89.82 39.06 89.92 39.16 ;
      RECT 89.82 39.27 89.92 39.37 ;
      RECT 89.82 39.48 89.92 39.58 ;
      RECT 89.82 39.69 89.92 39.79 ;
      RECT 89.61 39.06 89.71 39.16 ;
      RECT 89.61 39.27 89.71 39.37 ;
      RECT 89.61 39.48 89.71 39.58 ;
      RECT 89.61 39.69 89.71 39.79 ;
      RECT 89.4 39.06 89.5 39.16 ;
      RECT 89.4 39.27 89.5 39.37 ;
      RECT 89.4 39.48 89.5 39.58 ;
      RECT 89.4 39.69 89.5 39.79 ;
      RECT 82.36 0.1 82.46 0.2 ;
      RECT 82.36 0.3 82.46 0.4 ;
      RECT 82.12 0.1 82.22 0.2 ;
      RECT 82.12 0.3 82.22 0.4 ;
      RECT 81.1 39.15 81.2 39.25 ;
      RECT 81.1 39.35 81.2 39.45 ;
      RECT 81.1 39.55 81.2 39.65 ;
      RECT 81.1 39.75 81.2 39.85 ;
      RECT 80.86 39.15 80.96 39.25 ;
      RECT 80.86 39.35 80.96 39.45 ;
      RECT 80.86 39.55 80.96 39.65 ;
      RECT 80.86 39.75 80.96 39.85 ;
      RECT 63.63 39.055 63.73 39.155 ;
      RECT 63.63 39.265 63.73 39.365 ;
      RECT 63.63 39.475 63.73 39.575 ;
      RECT 63.63 39.685 63.73 39.785 ;
      RECT 63.42 39.055 63.52 39.155 ;
      RECT 63.42 39.265 63.52 39.365 ;
      RECT 63.42 39.475 63.52 39.575 ;
      RECT 63.42 39.685 63.52 39.785 ;
      RECT 63.21 39.055 63.31 39.155 ;
      RECT 63.21 39.265 63.31 39.365 ;
      RECT 63.21 39.475 63.31 39.575 ;
      RECT 63.21 39.685 63.31 39.785 ;
      RECT 63 39.055 63.1 39.155 ;
      RECT 63 39.265 63.1 39.365 ;
      RECT 63 39.475 63.1 39.575 ;
      RECT 63 39.685 63.1 39.785 ;
      RECT 62.79 39.055 62.89 39.155 ;
      RECT 62.79 39.265 62.89 39.365 ;
      RECT 62.79 39.475 62.89 39.575 ;
      RECT 62.79 39.685 62.89 39.785 ;
      RECT 62.58 39.055 62.68 39.155 ;
      RECT 62.58 39.265 62.68 39.365 ;
      RECT 62.58 39.475 62.68 39.575 ;
      RECT 62.58 39.685 62.68 39.785 ;
      RECT 58.915 39.06 59.015 39.16 ;
      RECT 58.915 39.27 59.015 39.37 ;
      RECT 58.915 39.48 59.015 39.58 ;
      RECT 58.915 39.69 59.015 39.79 ;
      RECT 58.705 39.06 58.805 39.16 ;
      RECT 58.705 39.27 58.805 39.37 ;
      RECT 58.705 39.48 58.805 39.58 ;
      RECT 58.705 39.69 58.805 39.79 ;
      RECT 58.495 39.06 58.595 39.16 ;
      RECT 58.495 39.27 58.595 39.37 ;
      RECT 58.495 39.48 58.595 39.58 ;
      RECT 58.495 39.69 58.595 39.79 ;
    LAYER ME3 ;
      RECT 88.19 35.59 89.19 37.74 ;
      RECT 81.45 35.59 82.55 37.74 ;
      RECT 57.86 35.59 58.26 37.8 ;
    LAYER ME3 SPACING 0.1 ;
      RECT 57.86 2.83 58.26 37.8 ;
      RECT 88.19 2.83 89.19 37.74 ;
      RECT 81.45 2.83 82.55 37.74 ;
      RECT 2.18 2.83 99.82 37.72 ;
      RECT 91.66 0 92.16 0.5 ;
      RECT 82.04 0 82.54 0.5 ;
    LAYER VI3 SPACING 0.1 ;
      RECT 1 1 101 38.9 ;
      RECT 91.98 0.1 92.08 0.2 ;
      RECT 91.98 0.3 92.08 0.4 ;
      RECT 91.74 0.1 91.84 0.2 ;
      RECT 91.74 0.3 91.84 0.4 ;
      RECT 82.36 0.1 82.46 0.2 ;
      RECT 82.36 0.3 82.46 0.4 ;
      RECT 82.12 0.1 82.22 0.2 ;
      RECT 82.12 0.3 82.22 0.4 ;
    LAYER ME4 SPACING 0.1 ;
      RECT 4.18 5.39 97.82 35.41 ;
      RECT 91.66 0 92.16 0.5 ;
      RECT 82.04 0 82.54 0.5 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END OSC_RINGTOPV1_NOVAR

END LIBRARY
