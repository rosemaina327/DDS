/**

This Module instantiates the analog physical components

*/
