/*

This module is the physical variant of the ADC, basically the same as the SPICE adc_analog module
*/
