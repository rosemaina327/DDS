module adc_analog (

    input wire VDD,
    input wire GND,

    input real VIN,
    input real VREF,

    output wire compout,
    input wire [7:0] vdac



);


endmodule
