/**
    Add the code for your adc_digital module here (SAR version)

*/
