module adc_analog (

    input wire VDD,
    input wire GND,

    input real VIN,
    input real VREF,

    input wire [7:0] vdac,

    output wire compout

);


endmodule
