`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AD42M2RA ( CO, ICO, S, A, B, C, D, ICI );
   input A, B, C, D, ICI;
   output CO, ICO, S;

    xor (tmp1, A, B, C);
    and (ts1,   D, tmp1);
    and (ts2, ICI, tmp1);
    and (ts3,   D,  ICI);
    or (CO, ts1, ts2, ts3);

    xor (tmp2, A, B);
    and (ts4,  tmp2, C);
    and (ts5,  A, B);
    or  (ICO, ts4, ts5);

     xor  (S, A, B, C, D, ICI);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc A --> ICO
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (A => ICO) = (0.0, 0.0);
    ifnone
        (A => ICO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (B => CO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (B => CO) = (0.0, 0.0);
    ifnone
        (B => CO) = (0.0, 0.0);

    // arc B --> ICO
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (B => ICO) = (0.0, 0.0);
    ifnone
        (B => ICO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc C --> CO
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1)
        (C => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0)
        (C => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
        (C => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
        (C => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
        (C => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
        (C => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1)
        (C => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0)
        (C => CO) = (0.0, 0.0);
    ifnone
        (C => CO) = (0.0, 0.0);

    // arc C --> ICO
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1)
        (C => ICO) = (0.0, 0.0);
    ifnone
        (C => ICO) = (0.0, 0.0);

    // arc C --> S
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    ifnone
        (C => S) = (0.0, 0.0);

    // arc D --> CO
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1)
        (D => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0)
        (D => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0)
        (D => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1)
        (D => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0)
        (D => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1)
        (D => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1)
        (D => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0)
        (D => CO) = (0.0, 0.0);
    ifnone
        (D => CO) = (0.0, 0.0);

    // arc D --> S
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    ifnone
        (D => S) = (0.0, 0.0);

    // arc ICI --> CO
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0)
        (ICI => CO) = (0.0, 0.0);
    ifnone
        (ICI => CO) = (0.0, 0.0);

    // arc ICI --> S
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    ifnone
        (ICI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AD42M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AD42M4RA ( CO, ICO, S, A, B, C, D, ICI );
   input A, B, C, D, ICI;
   output CO, ICO, S;

    xor (tmp1, A, B, C);
    and (ts1,   D, tmp1);
    and (ts2, ICI, tmp1);
    and (ts3,   D,  ICI);
    or (CO, ts1, ts2, ts3);

    xor (tmp2, A, B);
    and (ts4,  tmp2, C);
    and (ts5,  A, B);
    or  (ICO, ts4, ts5);

     xor  (S, A, B, C, D, ICI);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc A --> ICO
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (A => ICO) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (A => ICO) = (0.0, 0.0);
    ifnone
        (A => ICO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (B => CO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (B => CO) = (0.0, 0.0);
    ifnone
        (B => CO) = (0.0, 0.0);

    // arc B --> ICO
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (B => ICO) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (B => ICO) = (0.0, 0.0);
    ifnone
        (B => ICO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && ICI===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc C --> CO
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1)
        (C => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0)
        (C => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
        (C => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
        (C => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
        (C => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
        (C => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1)
        (C => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0)
        (C => CO) = (0.0, 0.0);
    ifnone
        (C => CO) = (0.0, 0.0);

    // arc C --> ICO
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
        (C => ICO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1)
        (C => ICO) = (0.0, 0.0);
    ifnone
        (C => ICO) = (0.0, 0.0);

    // arc C --> S
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b0 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b0)
        (C => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && ICI===1'b1)
        (C => S) = (0.0, 0.0);
    ifnone
        (C => S) = (0.0, 0.0);

    // arc D --> CO
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1)
        (D => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0)
        (D => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0)
        (D => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1)
        (D => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0)
        (D => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1)
        (D => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1)
        (D => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0)
        (D => CO) = (0.0, 0.0);
    ifnone
        (D => CO) = (0.0, 0.0);

    // arc D --> S
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b0 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b0)
        (D => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && ICI===1'b1)
        (D => S) = (0.0, 0.0);
    ifnone
        (D => S) = (0.0, 0.0);

    // arc ICI --> CO
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1)
        (ICI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0)
        (ICI => CO) = (0.0, 0.0);
    ifnone
        (ICI => CO) = (0.0, 0.0);

    // arc ICI --> S
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0)
        (ICI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b1)
        (ICI => S) = (0.0, 0.0);
    ifnone
        (ICI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AD42M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADCSCM2R ( CO0, CO1, A, B, NCI0, NCI1 );
   input A, B, NCI0, NCI1;
   output CO0, CO1;

         xor  (tmp1, A, B);
         and  (tmp2, A, B);
         not  (tmp3, NCI0);
         not  (tmp4, NCI1);
         and (ts1, tmp1,tmp3);
         or (CO0, ts1, tmp2);
         and (ts2, tmp1,tmp4);
         or (CO1, ts2, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    ifnone
        (A => CO0) = (0.0, 0.0);

    // arc A --> CO1
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    ifnone
        (A => CO1) = (0.0, 0.0);

    // arc B --> CO0
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    ifnone
        (B => CO0) = (0.0, 0.0);

    // arc B --> CO1
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    ifnone
        (B => CO1) = (0.0, 0.0);

    // arc NCI0 --> CO0
    if (A===1'b0 && B===1'b1 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    ifnone
        (NCI0 => CO0) = (0.0, 0.0);

    // arc NCI1 --> CO1
    if (A===1'b0 && B===1'b1 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    ifnone
        (NCI1 => CO1) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADCSCM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADCSCM4R ( CO0, CO1, A, B, NCI0, NCI1 );
   input A, B, NCI0, NCI1;
   output CO0, CO1;

         xor  (tmp1, A, B);
         and  (tmp2, A, B);
         not  (tmp3, NCI0);
         not  (tmp4, NCI1);
         and (ts1, tmp1,tmp3);
         or (CO0, ts1, tmp2);
         and (ts2, tmp1,tmp4);
         or (CO1, ts2, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    ifnone
        (A => CO0) = (0.0, 0.0);

    // arc A --> CO1
    if (B===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    ifnone
        (A => CO1) = (0.0, 0.0);

    // arc B --> CO0
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    ifnone
        (B => CO0) = (0.0, 0.0);

    // arc B --> CO1
    if (A===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    ifnone
        (B => CO1) = (0.0, 0.0);

    // arc NCI0 --> CO0
    if (A===1'b0 && B===1'b1 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    ifnone
        (NCI0 => CO0) = (0.0, 0.0);

    // arc NCI1 --> CO1
    if (A===1'b0 && B===1'b1 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    ifnone
        (NCI1 => CO1) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADCSCM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADCSIOM2R (A, B, CO0B, CO1B);
  input A, B;
  output CO0B, CO1B;

    nand SMC_I0(CO0B, A, B);

    not SMC_I1(A_bar, A);
    not SMC_I2(B_bar, B);
    and SMC_I3(CO1B, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    (A => CO0B) = (0.0, 0.0);

    // arc A --> CO1B
    (A => CO1B) = (0.0, 0.0);

    // arc B --> CO0B
    (B => CO0B) = (0.0, 0.0);

    // arc B --> CO1B
    (B => CO1B) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADCSIOM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADCSIOM4R (A, B, CO0B, CO1B);
  input A, B;
  output CO0B, CO1B;

    nand SMC_I0(CO0B, A, B);

    not SMC_I1(A_bar, A);
    not SMC_I2(B_bar, B);
    and SMC_I3(CO1B, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    (A => CO0B) = (0.0, 0.0);

    // arc A --> CO1B
    (A => CO1B) = (0.0, 0.0);

    // arc B --> CO0B
    (B => CO0B) = (0.0, 0.0);

    // arc B --> CO1B
    (B => CO1B) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADCSIOM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADCSOM2R ( CO0B, CO1B, A, B, CI0, CI1 );
   input A, B, CI0, CI1;
   output CO0B, CO1B;

       xor (tmp1, A, B);
       and (tmp2, A, B);
       and (ts1, tmp1, CI0);
       or (ts2, ts1, tmp2);
       not (CO0B, ts2);
       and (ts3, tmp1, CI1);
       or (ts4, ts3, tmp2);
       not (CO1B, ts4);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1)
        (A => CO0B) = (0.0, 0.0);
    ifnone
        (A => CO0B) = (0.0, 0.0);

    // arc A --> CO1B
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0)
        (A => CO1B) = (0.0, 0.0);
    ifnone
        (A => CO1B) = (0.0, 0.0);

    // arc B --> CO0B
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1)
        (B => CO0B) = (0.0, 0.0);
    ifnone
        (B => CO0B) = (0.0, 0.0);

    // arc B --> CO1B
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0)
        (B => CO1B) = (0.0, 0.0);
    ifnone
        (B => CO1B) = (0.0, 0.0);

    // arc CI0 --> CO0B
    if (A===1'b0 && B===1'b1 && CI1===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    ifnone
        (CI0 => CO0B) = (0.0, 0.0);

    // arc CI1 --> CO1B
    if (A===1'b0 && B===1'b1 && CI0===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    ifnone
        (CI1 => CO1B) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADCSOM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADCSOM4R ( CO0B, CO1B, A, B, CI0, CI1 );
   input A, B, CI0, CI1;
   output CO0B, CO1B;

       xor (tmp1, A, B);
       and (tmp2, A, B);
       and (ts1, tmp1, CI0);
       or (ts2, ts1, tmp2);
       not (CO0B, ts2);
       and (ts3, tmp1, CI1);
       or (ts4, ts3, tmp2);
       not (CO1B, ts4);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1)
        (A => CO0B) = (0.0, 0.0);
    ifnone
        (A => CO0B) = (0.0, 0.0);

    // arc A --> CO1B
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0)
        (A => CO1B) = (0.0, 0.0);
    ifnone
        (A => CO1B) = (0.0, 0.0);

    // arc B --> CO0B
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1)
        (B => CO0B) = (0.0, 0.0);
    ifnone
        (B => CO0B) = (0.0, 0.0);

    // arc B --> CO1B
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0)
        (B => CO1B) = (0.0, 0.0);
    ifnone
        (B => CO1B) = (0.0, 0.0);

    // arc CI0 --> CO0B
    if (A===1'b0 && B===1'b1 && CI1===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    ifnone
        (CI0 => CO0B) = (0.0, 0.0);

    // arc CI1 --> CO1B
    if (A===1'b0 && B===1'b1 && CI0===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    ifnone
        (CI1 => CO1B) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADCSOM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCGCM2RA ( CO, A, B, NCI );
   input A, B, NCI;
   output CO;

       xor (tmp1, A, B);
       and (tmp2, A, B);
       not (tmp3, NCI);
       and (ts1, tmp1, tmp3);
       or (CO, ts1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && NCI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && NCI===1'b1)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc B --> CO
    if (A===1'b0 && NCI===1'b0)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && NCI===1'b1)
        (B => CO) = (0.0, 0.0);
    ifnone
        (B => CO) = (0.0, 0.0);

    // arc NCI --> CO
    if (A===1'b0 && B===1'b1)
        (NCI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (NCI => CO) = (0.0, 0.0);
    ifnone
        (NCI => CO) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCGCM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCGCM4RA ( CO, A, B, NCI );
   input A, B, NCI;
   output CO;

       xor (tmp1, A, B);
       and (tmp2, A, B);
       not (tmp3, NCI);
       and (ts1, tmp1, tmp3);
       or (CO, ts1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && NCI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && NCI===1'b1)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc B --> CO
    if (A===1'b0 && NCI===1'b0)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && NCI===1'b1)
        (B => CO) = (0.0, 0.0);
    ifnone
        (B => CO) = (0.0, 0.0);

    // arc NCI --> CO
    if (A===1'b0 && B===1'b1)
        (NCI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (NCI => CO) = (0.0, 0.0);
    ifnone
        (NCI => CO) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCGCM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCGOM2RA ( COB, A, B, CI );
   input A, B, CI;
   output COB;

       xor (tmp1, A, B);
       and (tmp2, A, B);
       and (ts1, tmp1, CI);
       nor (COB, ts1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (B===1'b0 && CI===1'b1)
        (A => COB) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => COB) = (0.0, 0.0);
    ifnone
        (A => COB) = (0.0, 0.0);

    // arc B --> COB
    if (A===1'b0 && CI===1'b1)
        (B => COB) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => COB) = (0.0, 0.0);
    ifnone
        (B => COB) = (0.0, 0.0);

    // arc CI --> COB
    if (A===1'b0 && B===1'b1)
        (CI => COB) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => COB) = (0.0, 0.0);
    ifnone
        (CI => COB) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCGOM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCGOM4RA ( COB, A, B, CI );
   input A, B, CI;
   output COB;

       xor (tmp1, A, B);
       and (tmp2, A, B);
       and (ts1, tmp1, CI);
       nor (COB, ts1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (B===1'b0 && CI===1'b1)
        (A => COB) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => COB) = (0.0, 0.0);
    ifnone
        (A => COB) = (0.0, 0.0);

    // arc B --> COB
    if (A===1'b0 && CI===1'b1)
        (B => COB) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => COB) = (0.0, 0.0);
    ifnone
        (B => COB) = (0.0, 0.0);

    // arc CI --> COB
    if (A===1'b0 && B===1'b1)
        (CI => COB) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => COB) = (0.0, 0.0);
    ifnone
        (CI => COB) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCGOM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCM2RA ( CO, S, A, B, NCI );
   input A, B, NCI;
   output CO, S;

       xor (tmp1, A, B);
       and (tmp2, A, B);
       not (tmp3, NCI);
       and ( ts1, tmp1, tmp3);
       or ( CO, ts1, tmp2);
       xor ( S, tmp1, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && NCI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && NCI===1'b1)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && NCI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && NCI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && NCI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && NCI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    if (A===1'b0 && NCI===1'b0)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && NCI===1'b1)
        (B => CO) = (0.0, 0.0);
    ifnone
        (B => CO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && NCI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && NCI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && NCI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && NCI===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc NCI --> CO
    if (A===1'b0 && B===1'b1)
        (NCI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (NCI => CO) = (0.0, 0.0);
    ifnone
        (NCI => CO) = (0.0, 0.0);

    // arc NCI --> S
    if (A===1'b0 && B===1'b0)
        (NCI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (NCI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (NCI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (NCI => S) = (0.0, 0.0);
    ifnone
        (NCI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCM4RA ( CO, S, A, B, NCI );
   input A, B, NCI;
   output CO, S;

       xor (tmp1, A, B);
       and (tmp2, A, B);
       not (tmp3, NCI);
       and ( ts1, tmp1, tmp3);
       or ( CO, ts1, tmp2);
       xor ( S, tmp1, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && NCI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && NCI===1'b1)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && NCI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && NCI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && NCI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && NCI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    if (A===1'b0 && NCI===1'b0)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && NCI===1'b1)
        (B => CO) = (0.0, 0.0);
    ifnone
        (B => CO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && NCI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && NCI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && NCI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && NCI===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc NCI --> CO
    if (A===1'b0 && B===1'b1)
        (NCI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (NCI => CO) = (0.0, 0.0);
    ifnone
        (NCI => CO) = (0.0, 0.0);

    // arc NCI --> S
    if (A===1'b0 && B===1'b0)
        (NCI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (NCI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (NCI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (NCI => S) = (0.0, 0.0);
    ifnone
        (NCI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCSCM2RA ( CO0, CO1, S, A, B, CS, NCI0, NCI1 );
   input A, B, CS, NCI0, NCI1;
   output CO0, CO1, S;

      xor (tmp1, A, B);
      and (tmp2, A, B);
      not (tmp3, NCI0);
      not (tmp4, NCI1);
      not (tmp5, CS);
      and (ts1, tmp1, tmp3);
      or (CO0, ts1, tmp2);
      and (ts2, tmp1, tmp4);
      or (CO1, ts2, tmp2);
      xor (ts3, tmp1, tmp3);
      and (ts4, ts3, tmp5);
      xor (ts5, tmp1, tmp4);
      and (ts6, ts5, CS);
      or (S, ts4, ts6);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    ifnone
        (A => CO0) = (0.0, 0.0);

    // arc A --> CO1
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    ifnone
        (A => CO1) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO0
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    ifnone
        (B => CO0) = (0.0, 0.0);

    // arc B --> CO1
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    ifnone
        (B => CO1) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (CS => S) = (0.0, 0.0);
    ifnone
        (CS => S) = (0.0, 0.0);

    // arc NCI0 --> CO0
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    ifnone
        (NCI0 => CO0) = (0.0, 0.0);

    // arc NCI0 --> S
    if (A===1'b0 && B===1'b0 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => S) = (0.0, 0.0);
    ifnone
        (NCI0 => S) = (0.0, 0.0);

    // arc NCI1 --> CO1
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    ifnone
        (NCI1 => CO1) = (0.0, 0.0);

    // arc NCI1 --> S
    if (A===1'b0 && B===1'b0 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => S) = (0.0, 0.0);
    ifnone
        (NCI1 => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSCM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCSCM4RA ( CO0, CO1, S, A, B, CS, NCI0, NCI1 );
   input A, B, CS, NCI0, NCI1;
   output CO0, CO1, S;

      xor (tmp1, A, B);
      and (tmp2, A, B);
      not (tmp3, NCI0);
      not (tmp4, NCI1);
      not (tmp5, CS);
      and (ts1, tmp1, tmp3);
      or (CO0, ts1, tmp2);
      and (ts2, tmp1, tmp4);
      or (CO1, ts2, tmp2);
      xor (ts3, tmp1, tmp3);
      and (ts4, ts3, tmp5);
      xor (ts5, tmp1, tmp4);
      and (ts6, ts5, CS);
      or (S, ts4, ts6);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO0) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO0) = (0.0, 0.0);
    ifnone
        (A => CO0) = (0.0, 0.0);

    // arc A --> CO1
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => CO1) = (0.0, 0.0);
    ifnone
        (A => CO1) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO0
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO0) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO0) = (0.0, 0.0);
    ifnone
        (B => CO0) = (0.0, 0.0);

    // arc B --> CO1
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => CO1) = (0.0, 0.0);
    ifnone
        (B => CO1) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0 && NCI0===1'b1 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1 && NCI0===1'b1 && NCI1===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b0 && NCI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && NCI0===1'b1 && NCI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b0 && NCI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && NCI0===1'b1 && NCI1===1'b0)
        (CS => S) = (0.0, 0.0);
    ifnone
        (CS => S) = (0.0, 0.0);

    // arc NCI0 --> CO0
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b0)
        (NCI0 => CO0) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI1===1'b1)
        (NCI0 => CO0) = (0.0, 0.0);
    ifnone
        (NCI0 => CO0) = (0.0, 0.0);

    // arc NCI0 --> S
    if (A===1'b0 && B===1'b0 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CS===1'b0 && NCI1===1'b0)
        (NCI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CS===1'b0 && NCI1===1'b1)
        (NCI0 => S) = (0.0, 0.0);
    ifnone
        (NCI0 => S) = (0.0, 0.0);

    // arc NCI1 --> CO1
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b0 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b0 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => CO1) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => CO1) = (0.0, 0.0);
    ifnone
        (NCI1 => CO1) = (0.0, 0.0);

    // arc NCI1 --> S
    if (A===1'b0 && B===1'b0 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CS===1'b1 && NCI0===1'b0)
        (NCI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CS===1'b1 && NCI0===1'b1)
        (NCI1 => S) = (0.0, 0.0);
    ifnone
        (NCI1 => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSCM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCSIOM2R (A, B, CS, CO0B, CO1B, S);
  input A, B, CS;
  output CO0B, CO1B, S;

    nand SMC_I0(CO0B, A, B);

    not SMC_I1(A_bar, A);
    not SMC_I2(B_bar, B);
    and SMC_I3(CO1B, A_bar, B_bar);

    xor SMC_I4(S, A, B, CS);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (B===1'b1 && CS===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1)
        (A => CO0B) = (0.0, 0.0);
    ifnone
        (A => CO0B) = (0.0, 0.0);

    // arc A --> CO1B
    if (B===1'b0 && CS===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1)
        (A => CO1B) = (0.0, 0.0);
    ifnone
        (A => CO1B) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO0B
    if (A===1'b1 && CS===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (B => CO0B) = (0.0, 0.0);
    ifnone
        (B => CO0B) = (0.0, 0.0);

    // arc B --> CO1B
    if (A===1'b0 && CS===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1)
        (B => CO1B) = (0.0, 0.0);
    ifnone
        (B => CO1B) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (CS => S) = (0.0, 0.0);
    ifnone
        (CS => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSIOM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCSIOM4R (A, B, CS, CO0B, CO1B, S);
  input A, B, CS;
  output CO0B, CO1B, S;

    nand SMC_I0(CO0B, A, B);

    not SMC_I1(A_bar, A);
    not SMC_I2(B_bar, B);
    and SMC_I3(CO1B, A_bar, B_bar);

    xor SMC_I4(S, A, B, CS);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (B===1'b1 && CS===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1)
        (A => CO0B) = (0.0, 0.0);
    ifnone
        (A => CO0B) = (0.0, 0.0);

    // arc A --> CO1B
    if (B===1'b0 && CS===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1)
        (A => CO1B) = (0.0, 0.0);
    ifnone
        (A => CO1B) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO0B
    if (A===1'b1 && CS===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (B => CO0B) = (0.0, 0.0);
    ifnone
        (B => CO0B) = (0.0, 0.0);

    // arc B --> CO1B
    if (A===1'b0 && CS===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1)
        (B => CO1B) = (0.0, 0.0);
    ifnone
        (B => CO1B) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (CS => S) = (0.0, 0.0);
    ifnone
        (CS => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSIOM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCSOM2RA ( CO0B, CO1B, S, A, B, CI0, CI1, CS );
   input A, B, CI0, CI1, CS;
   output CO0B, CO1B, S;

     xor (tmp1, A, B);
     and (tmp2, A, B);
     not (tmp3, CS);
     and (ts1, tmp1, CI0);
     or (ts2, ts1, tmp2);
     not (CO0B, ts2);
     and (ts3, tmp1, CI1);
     or (ts4, ts3, tmp2);
     not (CO1B, ts4);
     xor (ts5, tmp1, CI0);
     and (ts6, ts5 , tmp3);
     xor (ts7, tmp1, CI1);
     and (ts8, ts7, CS);
     or (S, ts6, ts8);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (A => CO0B) = (0.0, 0.0);
    ifnone
        (A => CO0B) = (0.0, 0.0);

    // arc A --> CO1B
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (A => CO1B) = (0.0, 0.0);
    ifnone
        (A => CO1B) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO0B
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (B => CO0B) = (0.0, 0.0);
    ifnone
        (B => CO0B) = (0.0, 0.0);

    // arc B --> CO1B
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (B => CO1B) = (0.0, 0.0);
    ifnone
        (B => CO1B) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CI0 --> CO0B
    if (A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    ifnone
        (CI0 => CO0B) = (0.0, 0.0);

    // arc CI0 --> S
    if (A===1'b0 && B===1'b0 && CI1===1'b0 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && CI1===1'b1 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI1===1'b0 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI1===1'b1 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    ifnone
        (CI0 => S) = (0.0, 0.0);

    // arc CI1 --> CO1B
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    ifnone
        (CI1 => CO1B) = (0.0, 0.0);

    // arc CI1 --> S
    if (A===1'b0 && B===1'b0 && CI0===1'b0 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && CI0===1'b1 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b0 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b1 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    ifnone
        (CI1 => S) = (0.0, 0.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0 && CI0===1'b0 && CI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && CI0===1'b1 && CI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b0 && CI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b1 && CI1===1'b0)
        (CS => S) = (0.0, 0.0);
    ifnone
        (CS => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSOM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFCSOM4RA ( CO0B, CO1B, S, A, B, CI0, CI1, CS );
   input A, B, CI0, CI1, CS;
   output CO0B, CO1B, S;

     xor (tmp1, A, B);
     and (tmp2, A, B);
     not (tmp3, CS);
     and (ts1, tmp1, CI0);
     or (ts2, ts1, tmp2);
     not (CO0B, ts2);
     and (ts3, tmp1, CI1);
     or (ts4, ts3, tmp2);
     not (CO1B, ts4);
     xor (ts5, tmp1, CI0);
     and (ts6, ts5 , tmp3);
     xor (ts7, tmp1, CI1);
     and (ts8, ts7, CS);
     or (S, ts6, ts8);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO0B
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (A => CO0B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (A => CO0B) = (0.0, 0.0);
    ifnone
        (A => CO0B) = (0.0, 0.0);

    // arc A --> CO1B
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (A => CO1B) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (A => CO1B) = (0.0, 0.0);
    ifnone
        (A => CO1B) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO0B
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (B => CO0B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (B => CO0B) = (0.0, 0.0);
    ifnone
        (B => CO0B) = (0.0, 0.0);

    // arc B --> CO1B
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (B => CO1B) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (B => CO1B) = (0.0, 0.0);
    ifnone
        (B => CO1B) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b0 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b0 && CI1===1'b1 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b0 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI0===1'b1 && CI1===1'b1 && CS===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CI0 --> CO0B
    if (A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b0)
        (CI0 => CO0B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b1)
        (CI0 => CO0B) = (0.0, 0.0);
    ifnone
        (CI0 => CO0B) = (0.0, 0.0);

    // arc CI0 --> S
    if (A===1'b0 && B===1'b0 && CI1===1'b0 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && CI1===1'b1 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b0 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI1===1'b1 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b0 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI1===1'b1 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI1===1'b0 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI1===1'b1 && CS===1'b0)
        (CI0 => S) = (0.0, 0.0);
    ifnone
        (CI0 => S) = (0.0, 0.0);

    // arc CI1 --> CO1B
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b0)
        (CI1 => CO1B) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b1)
        (CI1 => CO1B) = (0.0, 0.0);
    ifnone
        (CI1 => CO1B) = (0.0, 0.0);

    // arc CI1 --> S
    if (A===1'b0 && B===1'b0 && CI0===1'b0 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && CI0===1'b1 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b0 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b1 && CS===1'b1)
        (CI1 => S) = (0.0, 0.0);
    ifnone
        (CI1 => S) = (0.0, 0.0);

    // arc CS --> S
    if (A===1'b0 && B===1'b0 && CI0===1'b0 && CI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && CI0===1'b1 && CI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b0 && CI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && CI0===1'b1 && CI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b0 && CI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && CI0===1'b1 && CI1===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b0 && CI1===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && CI0===1'b1 && CI1===1'b0)
        (CS => S) = (0.0, 0.0);
    ifnone
        (CS => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFCSOM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFM0RA ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;

      xor (tmp1, A, B);
      and (tmp2, A, B);
      and ( ts1, tmp1, CI);
      or ( CO, ts1, tmp2);
      xor ( S, A, B, CI);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => CO) = (0.0, 0.0);
    ifnone
        (B => CO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1)
        (CI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => CO) = (0.0, 0.0);
    ifnone
        (CI => CO) = (0.0, 0.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    ifnone
        (CI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFM0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFM1RA ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;

      xor (tmp1, A, B);
      and (tmp2, A, B);
      and ( ts1, tmp1, CI);
      or ( CO, ts1, tmp2);
      xor ( S, A, B, CI);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => CO) = (0.0, 0.0);
    ifnone
        (B => CO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1)
        (CI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => CO) = (0.0, 0.0);
    ifnone
        (CI => CO) = (0.0, 0.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    ifnone
        (CI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFM2RA ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;

      xor (tmp1, A, B);
      and (tmp2, A, B);
      and ( ts1, tmp1, CI);
      or ( CO, ts1, tmp2);
      xor ( S, A, B, CI);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => CO) = (0.0, 0.0);
    ifnone
        (B => CO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1)
        (CI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => CO) = (0.0, 0.0);
    ifnone
        (CI => CO) = (0.0, 0.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    ifnone
        (CI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFM4RA ( CO, S, A, B, CI );
   input A, B, CI;
   output CO, S;

      xor (tmp1, A, B);
      and (tmp2, A, B);
      and ( ts1, tmp1, CI);
      or ( CO, ts1, tmp2);
      xor ( S, A, B, CI);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (B===1'b0 && CI===1'b1)
        (A => CO) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    if (A===1'b0 && CI===1'b1)
        (B => CO) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => CO) = (0.0, 0.0);
    ifnone
        (B => CO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CI --> CO
    if (A===1'b0 && B===1'b1)
        (CI => CO) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => CO) = (0.0, 0.0);
    ifnone
        (CI => CO) = (0.0, 0.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    ifnone
        (CI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFOM2RA ( COB, S, A, B, CI );
   input A, B, CI;
   output COB, S;

      xor (tmp1, A, B);
      and (tmp2, A, B);
      and (ts1, tmp1, CI);
      or (ts2, ts1, tmp2);
      not (COB, ts2);
      xor (S, tmp1, CI);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (B===1'b0 && CI===1'b1)
        (A => COB) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => COB) = (0.0, 0.0);
    ifnone
        (A => COB) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> COB
    if (A===1'b0 && CI===1'b1)
        (B => COB) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => COB) = (0.0, 0.0);
    ifnone
        (B => COB) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CI --> COB
    if (A===1'b0 && B===1'b1)
        (CI => COB) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => COB) = (0.0, 0.0);
    ifnone
        (CI => COB) = (0.0, 0.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    ifnone
        (CI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFOM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADFOM4RA ( COB, S, A, B, CI );
   input A, B, CI;
   output COB, S;

      xor (tmp1, A, B);
      and (tmp2, A, B);
      and (ts1, tmp1, CI);
      or (ts2, ts1, tmp2);
      not (COB, ts2);
      xor (S, tmp1, CI);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (B===1'b0 && CI===1'b1)
        (A => COB) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => COB) = (0.0, 0.0);
    ifnone
        (A => COB) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b0 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1 && CI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> COB
    if (A===1'b0 && CI===1'b1)
        (B => COB) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => COB) = (0.0, 0.0);
    ifnone
        (B => COB) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b0 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);

    // arc CI --> COB
    if (A===1'b0 && B===1'b1)
        (CI => COB) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => COB) = (0.0, 0.0);
    ifnone
        (CI => COB) = (0.0, 0.0);

    // arc CI --> S
    if (A===1'b0 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (CI => S) = (0.0, 0.0);
    ifnone
        (CI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADFOM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCM2R (A, NCI, CO, S);
  input A, NCI;
  output CO, S;

    not SMC_I0(NCI_bar, NCI);
    and SMC_I1(CO, A, NCI_bar);

    xnor SMC_I2(S, A, NCI);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (NCI===1'b0)
        (A => S) = (0.0, 0.0);
    if (NCI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc NCI --> CO
    (NCI => CO) = (0.0, 0.0);

    // arc NCI --> S
    if (A===1'b0)
        (NCI => S) = (0.0, 0.0);
    if (A===1'b1)
        (NCI => S) = (0.0, 0.0);
    ifnone
        (NCI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHCM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCM4R (A, NCI, CO, S);
  input A, NCI;
  output CO, S;

    not SMC_I0(NCI_bar, NCI);
    and SMC_I1(CO, A, NCI_bar);

    xnor SMC_I2(S, A, NCI);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (NCI===1'b0)
        (A => S) = (0.0, 0.0);
    if (NCI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc NCI --> CO
    (NCI => CO) = (0.0, 0.0);

    // arc NCI --> S
    if (A===1'b0)
        (NCI => S) = (0.0, 0.0);
    if (A===1'b1)
        (NCI => S) = (0.0, 0.0);
    ifnone
        (NCI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHCM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCSCM2R (A, CS, NCI, CO, S);
  input A, CS, NCI;
  output CO, S;

    not SMC_I0(NCI_bar, NCI);
    and SMC_I1(CO, A, NCI_bar);

    not SMC_I2(A_bar, A);
    and SMC_I3(OUT0, A_bar, CS, NCI_bar);
    not SMC_I4(CS_bar, CS);
    and SMC_I5(OUT1, A, CS_bar);
    and SMC_I6(OUT2, A, NCI);
    or SMC_I7(S, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (CS===1'b0 && NCI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (CS===1'b1 && NCI===1'b0)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (CS===1'b0 && NCI===1'b0)
        (A => S) = (0.0, 0.0);
    if (CS===1'b0 && NCI===1'b1)
        (A => S) = (0.0, 0.0);
    if (CS===1'b1 && NCI===1'b0)
        (A => S) = (0.0, 0.0);
    if (CS===1'b1 && NCI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc CS --> S
    if (A===1'b0 && NCI===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && NCI===1'b0)
        (CS => S) = (0.0, 0.0);
    ifnone
        (CS => S) = (0.0, 0.0);

    // arc NCI --> CO
    if (A===1'b1 && CS===1'b0)
        (NCI => CO) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (NCI => CO) = (0.0, 0.0);
    ifnone
        (NCI => CO) = (0.0, 0.0);

    // arc NCI --> S
    if (A===1'b0 && CS===1'b1)
        (NCI => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (NCI => S) = (0.0, 0.0);
    ifnone
        (NCI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHCSCM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCSCM4R (A, CS, NCI, CO, S);
  input A, CS, NCI;
  output CO, S;

    not SMC_I0(NCI_bar, NCI);
    and SMC_I1(CO, A, NCI_bar);

    not SMC_I2(A_bar, A);
    and SMC_I3(OUT0, A_bar, CS, NCI_bar);
    not SMC_I4(CS_bar, CS);
    and SMC_I5(OUT1, A, CS_bar);
    and SMC_I6(OUT2, A, NCI);
    or SMC_I7(S, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    if (CS===1'b0 && NCI===1'b0)
        (A => CO) = (0.0, 0.0);
    if (CS===1'b1 && NCI===1'b0)
        (A => CO) = (0.0, 0.0);
    ifnone
        (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (CS===1'b0 && NCI===1'b0)
        (A => S) = (0.0, 0.0);
    if (CS===1'b0 && NCI===1'b1)
        (A => S) = (0.0, 0.0);
    if (CS===1'b1 && NCI===1'b0)
        (A => S) = (0.0, 0.0);
    if (CS===1'b1 && NCI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc CS --> S
    if (A===1'b0 && NCI===1'b0)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && NCI===1'b0)
        (CS => S) = (0.0, 0.0);
    ifnone
        (CS => S) = (0.0, 0.0);

    // arc NCI --> CO
    if (A===1'b1 && CS===1'b0)
        (NCI => CO) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (NCI => CO) = (0.0, 0.0);
    ifnone
        (NCI => CO) = (0.0, 0.0);

    // arc NCI --> S
    if (A===1'b0 && CS===1'b1)
        (NCI => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (NCI => S) = (0.0, 0.0);
    ifnone
        (NCI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHCSCM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCSOM2R (A, CI, CS, COB, S);
  input A, CI, CS;
  output COB, S;

    nand SMC_I0(COB, A, CI);

    not SMC_I1(CS_bar, CS);
    and SMC_I2(OUT0, A, CS_bar);
    not SMC_I3(CI_bar, CI);
    and SMC_I4(OUT1, A, CI_bar);
    not SMC_I5(A_bar, A);
    and SMC_I6(OUT2, A_bar, CI, CS);
    or SMC_I7(S, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (CI===1'b1 && CS===1'b0)
        (A => COB) = (0.0, 0.0);
    if (CI===1'b1 && CS===1'b1)
        (A => COB) = (0.0, 0.0);
    ifnone
        (A => COB) = (0.0, 0.0);

    // arc A --> S
    if (CI===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (CI===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (CI===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (CI===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc CI --> COB
    if (A===1'b1 && CS===1'b0)
        (CI => COB) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (CI => COB) = (0.0, 0.0);
    ifnone
        (CI => COB) = (0.0, 0.0);

    // arc CI --> S
    if (A===1'b0 && CS===1'b1)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (CI => S) = (0.0, 0.0);
    ifnone
        (CI => S) = (0.0, 0.0);

    // arc CS --> S
    if (A===1'b0 && CI===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b1)
        (CS => S) = (0.0, 0.0);
    ifnone
        (CS => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHCSOM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHCSOM4R (A, CI, CS, COB, S);
  input A, CI, CS;
  output COB, S;

    nand SMC_I0(COB, A, CI);

    not SMC_I1(CS_bar, CS);
    and SMC_I2(OUT0, A, CS_bar);
    not SMC_I3(CI_bar, CI);
    and SMC_I4(OUT1, A, CI_bar);
    not SMC_I5(A_bar, A);
    and SMC_I6(OUT2, A_bar, CI, CS);
    or SMC_I7(S, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    if (CI===1'b1 && CS===1'b0)
        (A => COB) = (0.0, 0.0);
    if (CI===1'b1 && CS===1'b1)
        (A => COB) = (0.0, 0.0);
    ifnone
        (A => COB) = (0.0, 0.0);

    // arc A --> S
    if (CI===1'b0 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (CI===1'b0 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    if (CI===1'b1 && CS===1'b0)
        (A => S) = (0.0, 0.0);
    if (CI===1'b1 && CS===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc CI --> COB
    if (A===1'b1 && CS===1'b0)
        (CI => COB) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (CI => COB) = (0.0, 0.0);
    ifnone
        (CI => COB) = (0.0, 0.0);

    // arc CI --> S
    if (A===1'b0 && CS===1'b1)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1 && CS===1'b1)
        (CI => S) = (0.0, 0.0);
    ifnone
        (CI => S) = (0.0, 0.0);

    // arc CS --> S
    if (A===1'b0 && CI===1'b1)
        (CS => S) = (0.0, 0.0);
    if (A===1'b1 && CI===1'b1)
        (CS => S) = (0.0, 0.0);
    ifnone
        (CS => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHCSOM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHM1RA (A, B, CO, S);
  input A, B;
  output CO, S;

    and SMC_I0(CO, A, B);

    xor SMC_I1(S, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    (B => CO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHM2RA (A, B, CO, S);
  input A, B;
  output CO, S;

    and SMC_I0(CO, A, B);

    xor SMC_I1(S, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    (B => CO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHM4RA (A, B, CO, S);
  input A, B;
  output CO, S;

    and SMC_I0(CO, A, B);

    xor SMC_I1(S, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    (B => CO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHM8RA (A, B, CO, S);
  input A, B;
  output CO, S;

    and SMC_I0(CO, A, B);

    xor SMC_I1(S, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> CO
    (A => CO) = (0.0, 0.0);

    // arc A --> S
    if (B===1'b0)
        (A => S) = (0.0, 0.0);
    if (B===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc B --> CO
    (B => CO) = (0.0, 0.0);

    // arc B --> S
    if (A===1'b0)
        (B => S) = (0.0, 0.0);
    if (A===1'b1)
        (B => S) = (0.0, 0.0);
    ifnone
        (B => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHOM2R (A, CI, COB, S);
  input A, CI;
  output COB, S;

    nand SMC_I0(COB, A, CI);

    xor SMC_I1(S, A, CI);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    (A => COB) = (0.0, 0.0);

    // arc A --> S
    if (CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (CI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc CI --> COB
    (CI => COB) = (0.0, 0.0);

    // arc CI --> S
    if (A===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1)
        (CI => S) = (0.0, 0.0);
    ifnone
        (CI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHOM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ADHOM4R (A, CI, COB, S);
  input A, CI;
  output COB, S;

    nand SMC_I0(COB, A, CI);

    xor SMC_I1(S, A, CI);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> COB
    (A => COB) = (0.0, 0.0);

    // arc A --> S
    if (CI===1'b0)
        (A => S) = (0.0, 0.0);
    if (CI===1'b1)
        (A => S) = (0.0, 0.0);
    ifnone
        (A => S) = (0.0, 0.0);

    // arc CI --> COB
    (CI => COB) = (0.0, 0.0);

    // arc CI --> S
    if (A===1'b0)
        (CI => S) = (0.0, 0.0);
    if (A===1'b1)
        (CI => S) = (0.0, 0.0);
    ifnone
        (CI => S) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ADHOM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M0R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN2M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M12RA (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN2M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M16RA (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN2M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M1R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN2M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M22RA (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN2M22RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M2R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN2M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M4R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN2M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M6R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN2M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN2M8R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN2M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN3M0R ( Z, A, B, C );
   input A, B, C;
   output Z;

    and (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN3M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN3M12RA ( Z, A, B, C );
   input A, B, C;
   output Z;

    and (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN3M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN3M16RA ( Z, A, B, C );
   input A, B, C;
   output Z;

    and (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN3M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN3M1R ( Z, A, B, C );
   input A, B, C;
   output Z;

    and (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN3M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN3M22RA ( Z, A, B, C );
   input A, B, C;
   output Z;

    and (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN3M22RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN3M2R ( Z, A, B, C );
   input A, B, C;
   output Z;

    and (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN3M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN3M4R ( Z, A, B, C );
   input A, B, C;
   output Z;

    and (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN3M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN3M6R ( Z, A, B, C );
   input A, B, C;
   output Z;

    and (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN3M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN3M8R ( Z, A, B, C );
   input A, B, C;
   output Z;

    and (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN3M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN4M0R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    and (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN4M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN4M12RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    and (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN4M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN4M16RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    and (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN4M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN4M1R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    and (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN4M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN4M2R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    and (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN4M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN4M4RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    and (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN4M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN4M6R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    and (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN4M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AN4M8RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    and (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AN4M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO211M1RA (A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, C);
    buf SMC_I2(OUT2, B);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO211M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO211M2RA (A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, C);
    buf SMC_I2(OUT2, B);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO211M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO211M4RA (A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, C);
    buf SMC_I2(OUT2, B);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO211M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO211M8RA (A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, C);
    buf SMC_I2(OUT2, B);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO211M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M0RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO21M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M12RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO21M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M1RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO21M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M2RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO21M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M4RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO21M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M6RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO21M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO21M8RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, A2);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO21M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO221M1RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      AO221_UDP5(Z, A1, A2, B1, B2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO221M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO221M2RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      AO221_UDP5(Z, A1, A2, B1, B2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO221M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO221M4RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      AO221_UDP5(Z, A1, A2, B1, B2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO221M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO221M8RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      AO221_UDP5(Z, A1, A2, B1, B2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO221M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO222M1RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      AO222_UDP6(Z, A1, A2, B1, B2, C1, C2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO222M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO222M2RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      AO222_UDP6(Z, A1, A2, B1, B2, C1, C2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO222M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO222M4RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      AO222_UDP6(Z, A1, A2, B1, B2, C1, C2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO222M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO222M8RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      AO222_UDP6(Z, A1, A2, B1, B2, C1, C2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO222M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22B10M0R ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;

    not (tmp1, NA2);
    and (tmp2, A1, tmp1);
    and (tmp3, B1, B2);
    or (Z, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && B2===1'b0 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && B2===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B2===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && B1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22B10M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22B10M1R ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;

    not (tmp1, NA2);
    and (tmp2, A1, tmp1);
    and (tmp3, B1, B2);
    or (Z, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && B2===1'b0 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && B2===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B2===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && B1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22B10M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22B10M2R ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;

    not (tmp1, NA2);
    and (tmp2, A1, tmp1);
    and (tmp3, B1, B2);
    or (Z, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && B2===1'b0 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && B2===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B2===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && B1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22B10M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22B10M4R ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;

    not (tmp1, NA2);
    and (tmp2, A1, tmp1);
    and (tmp3, B1, B2);
    or (Z, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && B2===1'b0 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && B2===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B2===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && B1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22B10M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22B10M8RA ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;

    not (tmp1, NA2);
    and (tmp2, A1, tmp1);
    and (tmp3, B1, B2);
    or (Z, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && B2===1'b0 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && B2===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B2===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && B1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22B10M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22B11M0R ( Z, A1, B1, NA2, NB2 );
   input A1, B1, NA2, NB2;
   output Z;

    not (tmp1, NA2);
    not (tmp2, NB2);
    and (ts1, A1, tmp1);
    and (ts2, B1, tmp2);
    or (Z, ts1, ts2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && NA2===1'b0 && NB2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA2===1'b0 && NB2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA2===1'b0 && NB2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && NA2===1'b0 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b1 && B1===1'b0 && NB2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NB2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NB2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);

    // arc NB2 --> Z
    if (A1===1'b0 && B1===1'b1 && NA2===1'b0)
        (NB2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && NA2===1'b1)
        (NB2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NA2===1'b1)
        (NB2 => Z) = (0.0, 0.0);
    ifnone
        (NB2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22B11M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22B11M1R ( Z, A1, B1, NA2, NB2 );
   input A1, B1, NA2, NB2;
   output Z;

    not (tmp1, NA2);
    not (tmp2, NB2);
    and (ts1, A1, tmp1);
    and (ts2, B1, tmp2);
    or (Z, ts1, ts2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && NA2===1'b0 && NB2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA2===1'b0 && NB2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA2===1'b0 && NB2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && NA2===1'b0 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b1 && B1===1'b0 && NB2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NB2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NB2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);

    // arc NB2 --> Z
    if (A1===1'b0 && B1===1'b1 && NA2===1'b0)
        (NB2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && NA2===1'b1)
        (NB2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NA2===1'b1)
        (NB2 => Z) = (0.0, 0.0);
    ifnone
        (NB2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22B11M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22B11M2R ( Z, A1, B1, NA2, NB2 );
   input A1, B1, NA2, NB2;
   output Z;

    not (tmp1, NA2);
    not (tmp2, NB2);
    and (ts1, A1, tmp1);
    and (ts2, B1, tmp2);
    or (Z, ts1, ts2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && NA2===1'b0 && NB2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA2===1'b0 && NB2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA2===1'b0 && NB2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && NA2===1'b0 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b1 && B1===1'b0 && NB2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NB2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NB2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);

    // arc NB2 --> Z
    if (A1===1'b0 && B1===1'b1 && NA2===1'b0)
        (NB2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && NA2===1'b1)
        (NB2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NA2===1'b1)
        (NB2 => Z) = (0.0, 0.0);
    ifnone
        (NB2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22B11M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22B11M4R ( Z, A1, B1, NA2, NB2 );
   input A1, B1, NA2, NB2;
   output Z;

    not (tmp1, NA2);
    not (tmp2, NB2);
    and (ts1, A1, tmp1);
    and (ts2, B1, tmp2);
    or (Z, ts1, ts2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && NA2===1'b0 && NB2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA2===1'b0 && NB2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA2===1'b0 && NB2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && NA2===1'b0 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b1 && B1===1'b0 && NB2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NB2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NB2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);

    // arc NB2 --> Z
    if (A1===1'b0 && B1===1'b1 && NA2===1'b0)
        (NB2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && NA2===1'b1)
        (NB2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NA2===1'b1)
        (NB2 => Z) = (0.0, 0.0);
    ifnone
        (NB2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22B11M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22B11M8RA ( Z, A1, B1, NA2, NB2 );
   input A1, B1, NA2, NB2;
   output Z;

    not (tmp1, NA2);
    not (tmp2, NB2);
    and (ts1, A1, tmp1);
    and (ts2, B1, tmp2);
    or (Z, ts1, ts2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && NA2===1'b0 && NB2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA2===1'b0 && NB2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA2===1'b0 && NB2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && NA2===1'b0 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1 && NB2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b1 && B1===1'b0 && NB2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NB2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NB2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);

    // arc NB2 --> Z
    if (A1===1'b0 && B1===1'b1 && NA2===1'b0)
        (NB2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && NA2===1'b1)
        (NB2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && NA2===1'b1)
        (NB2 => Z) = (0.0, 0.0);
    ifnone
        (NB2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22B11M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22M0RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

    and ( tmp1, A1, A2);
    and ( tmp2, B1, B2);
     or (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22M12RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

    and ( tmp1, A1, A2);
    and ( tmp2, B1, B2);
     or (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22M1RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

    and ( tmp1, A1, A2);
    and ( tmp2, B1, B2);
     or (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22M2R ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

    and ( tmp1, A1, A2);
    and ( tmp2, B1, B2);
     or (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22M4RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

    and ( tmp1, A1, A2);
    and ( tmp2, B1, B2);
     or (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22M6RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

    and ( tmp1, A1, A2);
    and ( tmp2, B1, B2);
     or (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO22M8RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

    and ( tmp1, A1, A2);
    and ( tmp2, B1, B2);
     or (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO22M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO31M1RA ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;
      AO31_UDP4(Z, A1, A2, A3, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO31M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO31M2RA ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;
      AO31_UDP4(Z, A1, A2, A3, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO31M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO31M4RA ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;
      AO31_UDP4(Z, A1, A2, A3, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO31M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO31M8RA ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;
      AO31_UDP4(Z, A1, A2, A3, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO31M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO32M1RA ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;
      AO32_UDP5(Z, A1, A2, A3, B1, B2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO32M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO32M2RA ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;
      AO32_UDP5(Z, A1, A2, A3, B1, B2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO32M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO32M4RA ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;
      AO32_UDP5(Z, A1, A2, A3, B1, B2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO32M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO32M8RA ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;
      AO32_UDP5(Z, A1, A2, A3, B1, B2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO32M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO33M1RA ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;
      AO33_UDP6(Z, A1, A2, A3, B1, B2, B3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO33M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO33M2RA ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;
      AO33_UDP6(Z, A1, A2, A3, B1, B2, B3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO33M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO33M4RA ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;
      AO33_UDP6(Z, A1, A2, A3, B1, B2, B3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO33M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AO33M8RA ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;
      AO33_UDP6(Z, A1, A2, A3, B1, B2, B3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AO33M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI211M0R ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI211M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI211M1R ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI211M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI211M2R ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI211M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI211M4R ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI211M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI211M6RA ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI211M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI211M8RA ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI211M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M0R (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M12RA (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M16RA (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M1R (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M2R (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M4R (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M6RA (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B01M8RA (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, NB);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B01M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M0R (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M12RA (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M16RA (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M1R (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M2R (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M4R (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M6RA (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B10M8RA (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A1_bar, B_bar);
    and SMC_I3(OUT1, B_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B10M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B20M0R (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(OUT0, B_bar, NA2);
    and SMC_I2(OUT1, B_bar, NA1);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B20M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B20M1R (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(OUT0, B_bar, NA2);
    and SMC_I2(OUT1, B_bar, NA1);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B20M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B20M2R (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(OUT0, B_bar, NA2);
    and SMC_I2(OUT1, B_bar, NA1);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B20M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B20M4R (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(OUT0, B_bar, NA2);
    and SMC_I2(OUT1, B_bar, NA1);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B20M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21B20M8RA (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(OUT0, B_bar, NA2);
    and SMC_I2(OUT1, B_bar, NA1);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21B20M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M0R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M12RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M16RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M1R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M2R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M3R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M4R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M6R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI21M8R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

     and (tmp1, A1, A2);
     nor (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI21M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI221M0R ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    nor (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI221M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI221M1R ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    nor (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI221M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI221M2R ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    nor (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI221M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI221M4R ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    nor (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI221M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI221M6RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    nor (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI221M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI221M8RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    nor (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI221M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI222M0RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    and (tmp3, C1, C2);
    nor (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI222M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI222M1RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    and (tmp3, C1, C2);
    nor (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI222M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI222M2R ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    and (tmp3, C1, C2);
    nor (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI222M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI222M4R ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    and (tmp3, C1, C2);
    nor (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI222M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI222M6RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    and (tmp3, C1, C2);
    nor (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI222M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI222M8RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

    and (tmp1, A1, A2);
    and (tmp2, B1, B2);
    and (tmp3, C1, C2);
    nor (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b1)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI222M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22B20M0R (B1, B2, NA1, NA2, Z);
  input B1, B2, NA1, NA2;
  output Z;

    not SMC_I0(B1_bar, B1);
    and SMC_I1(OUT0, B1_bar, NA1);
    not SMC_I2(B2_bar, B2);
    and SMC_I3(OUT1, B2_bar, NA1);
    and SMC_I4(OUT2, B1_bar, NA2);
    and SMC_I5(OUT3, B2_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    if (B2===1'b1 && NA1===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b1 && NA1===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b1 && NA1===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (B1===1'b1 && NA1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    if (B1===1'b0 && B2===1'b0 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    ifnone
        (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (B1===1'b0 && B2===1'b0 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22B20M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22B20M1R (B1, B2, NA1, NA2, Z);
  input B1, B2, NA1, NA2;
  output Z;

    not SMC_I0(B1_bar, B1);
    and SMC_I1(OUT0, B1_bar, NA1);
    not SMC_I2(B2_bar, B2);
    and SMC_I3(OUT1, B2_bar, NA1);
    and SMC_I4(OUT2, B1_bar, NA2);
    and SMC_I5(OUT3, B2_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    if (B2===1'b1 && NA1===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b1 && NA1===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b1 && NA1===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (B1===1'b1 && NA1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    if (B1===1'b0 && B2===1'b0 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    ifnone
        (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (B1===1'b0 && B2===1'b0 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22B20M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22B20M2R (B1, B2, NA1, NA2, Z);
  input B1, B2, NA1, NA2;
  output Z;

    not SMC_I0(B1_bar, B1);
    and SMC_I1(OUT0, B1_bar, NA1);
    not SMC_I2(B2_bar, B2);
    and SMC_I3(OUT1, B2_bar, NA1);
    and SMC_I4(OUT2, B1_bar, NA2);
    and SMC_I5(OUT3, B2_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    if (B2===1'b1 && NA1===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b1 && NA1===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b1 && NA1===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (B1===1'b1 && NA1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    if (B1===1'b0 && B2===1'b0 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    ifnone
        (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (B1===1'b0 && B2===1'b0 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22B20M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22B20M4R (B1, B2, NA1, NA2, Z);
  input B1, B2, NA1, NA2;
  output Z;

    not SMC_I0(B1_bar, B1);
    and SMC_I1(OUT0, B1_bar, NA1);
    not SMC_I2(B2_bar, B2);
    and SMC_I3(OUT1, B2_bar, NA1);
    and SMC_I4(OUT2, B1_bar, NA2);
    and SMC_I5(OUT3, B2_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    if (B2===1'b1 && NA1===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b1 && NA1===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b1 && NA1===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (B1===1'b1 && NA1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    if (B1===1'b0 && B2===1'b0 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    ifnone
        (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (B1===1'b0 && B2===1'b0 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22B20M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22B20M8RA (B1, B2, NA1, NA2, Z);
  input B1, B2, NA1, NA2;
  output Z;

    not SMC_I0(B1_bar, B1);
    and SMC_I1(OUT0, B1_bar, NA1);
    not SMC_I2(B2_bar, B2);
    and SMC_I3(OUT1, B2_bar, NA1);
    and SMC_I4(OUT2, B1_bar, NA2);
    and SMC_I5(OUT3, B2_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    if (B2===1'b1 && NA1===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b1 && NA1===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b1 && NA1===1'b1 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (B1===1'b1 && NA1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && NA1===1'b1 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    if (B1===1'b0 && B2===1'b0 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b0)
        (NA1 => Z) = (0.0, 0.0);
    ifnone
        (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (B1===1'b0 && B2===1'b0 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && B2===1'b1 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA1===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22B20M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M0R (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M12RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M16RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M1R (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M2R (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M4R (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M6RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI22M8RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B1_bar);
    not SMC_I5(B2_bar, B2);
    and SMC_I6(OUT2, A2_bar, B2_bar);
    and SMC_I7(OUT3, A1_bar, B2_bar);
    or SMC_I8(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI22M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M0R (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M12RA (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M1R (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M2R (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M4R (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M6RA (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI31M8RA (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    not SMC_I0(A3_bar, A3);
    not SMC_I1(B_bar, B);
    and SMC_I2(OUT0, A3_bar, B_bar);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A2_bar, B_bar);
    not SMC_I5(A1_bar, A1);
    and SMC_I6(OUT2, A1_bar, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI31M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M0R (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M12RA (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M1R (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M2R (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M4R (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M6RA (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI32M8RA (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B2_bar, B2);
    and SMC_I2(OUT0, A1_bar, B2_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B1_bar, B1);
    and SMC_I5(OUT1, A3_bar, B1_bar);
    and SMC_I6(OUT2, A1_bar, B1_bar);
    and SMC_I7(OUT3, A3_bar, B2_bar);
    not SMC_I8(A2_bar, A2);
    and SMC_I9(OUT4, A2_bar, B1_bar);
    and SMC_I10(OUT5, A2_bar, B2_bar);
    or SMC_I11(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI32M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI33M0R (A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B3_bar, B3);
    and SMC_I5(OUT1, A3_bar, B3_bar);
    and SMC_I6(OUT2, A1_bar, B3_bar);
    not SMC_I7(A2_bar, A2);
    and SMC_I8(OUT3, A2_bar, B1_bar);
    not SMC_I9(B2_bar, B2);
    and SMC_I10(OUT4, A3_bar, B2_bar);
    and SMC_I11(OUT5, A2_bar, B2_bar);
    and SMC_I12(OUT6, A2_bar, B3_bar);
    and SMC_I13(OUT7, A3_bar, B1_bar);
    and SMC_I14(OUT8, A1_bar, B2_bar);
    or SMC_I15(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I16(OUTSUB1, OUT8);
    or SMC_I17(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI33M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI33M1R (A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B3_bar, B3);
    and SMC_I5(OUT1, A3_bar, B3_bar);
    and SMC_I6(OUT2, A1_bar, B3_bar);
    not SMC_I7(A2_bar, A2);
    and SMC_I8(OUT3, A2_bar, B1_bar);
    not SMC_I9(B2_bar, B2);
    and SMC_I10(OUT4, A3_bar, B2_bar);
    and SMC_I11(OUT5, A2_bar, B2_bar);
    and SMC_I12(OUT6, A2_bar, B3_bar);
    and SMC_I13(OUT7, A3_bar, B1_bar);
    and SMC_I14(OUT8, A1_bar, B2_bar);
    or SMC_I15(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I16(OUTSUB1, OUT8);
    or SMC_I17(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI33M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI33M2R (A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B3_bar, B3);
    and SMC_I5(OUT1, A3_bar, B3_bar);
    and SMC_I6(OUT2, A1_bar, B3_bar);
    not SMC_I7(A2_bar, A2);
    and SMC_I8(OUT3, A2_bar, B1_bar);
    not SMC_I9(B2_bar, B2);
    and SMC_I10(OUT4, A3_bar, B2_bar);
    and SMC_I11(OUT5, A2_bar, B2_bar);
    and SMC_I12(OUT6, A2_bar, B3_bar);
    and SMC_I13(OUT7, A3_bar, B1_bar);
    and SMC_I14(OUT8, A1_bar, B2_bar);
    or SMC_I15(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I16(OUTSUB1, OUT8);
    or SMC_I17(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI33M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI33M4R (A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B3_bar, B3);
    and SMC_I5(OUT1, A3_bar, B3_bar);
    and SMC_I6(OUT2, A1_bar, B3_bar);
    not SMC_I7(A2_bar, A2);
    and SMC_I8(OUT3, A2_bar, B1_bar);
    not SMC_I9(B2_bar, B2);
    and SMC_I10(OUT4, A3_bar, B2_bar);
    and SMC_I11(OUT5, A2_bar, B2_bar);
    and SMC_I12(OUT6, A2_bar, B3_bar);
    and SMC_I13(OUT7, A3_bar, B1_bar);
    and SMC_I14(OUT8, A1_bar, B2_bar);
    or SMC_I15(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I16(OUTSUB1, OUT8);
    or SMC_I17(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI33M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module AOI33M8RA (A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(B1_bar, B1);
    and SMC_I2(OUT0, A1_bar, B1_bar);
    not SMC_I3(A3_bar, A3);
    not SMC_I4(B3_bar, B3);
    and SMC_I5(OUT1, A3_bar, B3_bar);
    and SMC_I6(OUT2, A1_bar, B3_bar);
    not SMC_I7(A2_bar, A2);
    and SMC_I8(OUT3, A2_bar, B1_bar);
    not SMC_I9(B2_bar, B2);
    and SMC_I10(OUT4, A3_bar, B2_bar);
    and SMC_I11(OUT5, A2_bar, B2_bar);
    and SMC_I12(OUT6, A2_bar, B3_bar);
    and SMC_I13(OUT7, A3_bar, B1_bar);
    and SMC_I14(OUT8, A1_bar, B2_bar);
    or SMC_I15(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I16(OUTSUB1, OUT8);
    or SMC_I17(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b1 && B3===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B3===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // AOI33M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEM2RA (M0, M1, M2, OA1, OA2, Z);
  input M0, M1, M2;
  output OA1, OA2, Z;

    and SMC_I0(OUT0, M0, M1);
    not SMC_I1(M2_bar, M2);
    buf SMC_I2(OUT1, M2_bar);
    or SMC_I3(OA1, OUT0, OUT1);

    not SMC_I4(M0_bar, M0);
    not SMC_I5(M1_bar, M1);
    and SMC_I6(OUT2, M0_bar, M1_bar);
    buf SMC_I7(OUT3, M2);
    or SMC_I8(OA2, OUT2, OUT3);

    xnor SMC_I9(Z, M0, M1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> OA1
    (M0 => OA1) = (0.0, 0.0);

    // arc M0 --> OA2
    (M0 => OA2) = (0.0, 0.0);

    // arc M0 --> Z
    if (M1===1'b0 && M2===1'b0)
        (M0 => Z) = (0.0, 0.0);
    if (M1===1'b0 && M2===1'b1)
        (M0 => Z) = (0.0, 0.0);
    if (M1===1'b1 && M2===1'b0)
        (M0 => Z) = (0.0, 0.0);
    if (M1===1'b1 && M2===1'b1)
        (M0 => Z) = (0.0, 0.0);
    ifnone
        (M0 => Z) = (0.0, 0.0);

    // arc M1 --> OA1
    (M1 => OA1) = (0.0, 0.0);

    // arc M1 --> OA2
    (M1 => OA2) = (0.0, 0.0);

    // arc M1 --> Z
    if (M0===1'b0 && M2===1'b0)
        (M1 => Z) = (0.0, 0.0);
    if (M0===1'b0 && M2===1'b1)
        (M1 => Z) = (0.0, 0.0);
    if (M0===1'b1 && M2===1'b0)
        (M1 => Z) = (0.0, 0.0);
    if (M0===1'b1 && M2===1'b1)
        (M1 => Z) = (0.0, 0.0);
    ifnone
        (M1 => Z) = (0.0, 0.0);

    // arc M2 --> OA1
    if (M0===1'b0 && M1===1'b0)
        (M2 => OA1) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1)
        (M2 => OA1) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0)
        (M2 => OA1) = (0.0, 0.0);
    ifnone
        (M2 => OA1) = (0.0, 0.0);

    // arc M2 --> OA2
    if (M0===1'b0 && M1===1'b1)
        (M2 => OA2) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0)
        (M2 => OA2) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1)
        (M2 => OA2) = (0.0, 0.0);
    ifnone
        (M2 => OA2) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BEM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEM4RA (M0, M1, M2, OA1, OA2, Z);
  input M0, M1, M2;
  output OA1, OA2, Z;

    and SMC_I0(OUT0, M0, M1);
    not SMC_I1(M2_bar, M2);
    buf SMC_I2(OUT1, M2_bar);
    or SMC_I3(OA1, OUT0, OUT1);

    not SMC_I4(M0_bar, M0);
    not SMC_I5(M1_bar, M1);
    and SMC_I6(OUT2, M0_bar, M1_bar);
    buf SMC_I7(OUT3, M2);
    or SMC_I8(OA2, OUT2, OUT3);

    xnor SMC_I9(Z, M0, M1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> OA1
    (M0 => OA1) = (0.0, 0.0);

    // arc M0 --> OA2
    (M0 => OA2) = (0.0, 0.0);

    // arc M0 --> Z
    if (M1===1'b0 && M2===1'b0)
        (M0 => Z) = (0.0, 0.0);
    if (M1===1'b0 && M2===1'b1)
        (M0 => Z) = (0.0, 0.0);
    if (M1===1'b1 && M2===1'b0)
        (M0 => Z) = (0.0, 0.0);
    if (M1===1'b1 && M2===1'b1)
        (M0 => Z) = (0.0, 0.0);
    ifnone
        (M0 => Z) = (0.0, 0.0);

    // arc M1 --> OA1
    (M1 => OA1) = (0.0, 0.0);

    // arc M1 --> OA2
    (M1 => OA2) = (0.0, 0.0);

    // arc M1 --> Z
    if (M0===1'b0 && M2===1'b0)
        (M1 => Z) = (0.0, 0.0);
    if (M0===1'b0 && M2===1'b1)
        (M1 => Z) = (0.0, 0.0);
    if (M0===1'b1 && M2===1'b0)
        (M1 => Z) = (0.0, 0.0);
    if (M0===1'b1 && M2===1'b1)
        (M1 => Z) = (0.0, 0.0);
    ifnone
        (M1 => Z) = (0.0, 0.0);

    // arc M2 --> OA1
    if (M0===1'b0 && M1===1'b0)
        (M2 => OA1) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1)
        (M2 => OA1) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0)
        (M2 => OA1) = (0.0, 0.0);
    ifnone
        (M2 => OA1) = (0.0, 0.0);

    // arc M2 --> OA2
    if (M0===1'b0 && M1===1'b1)
        (M2 => OA2) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0)
        (M2 => OA2) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1)
        (M2 => OA2) = (0.0, 0.0);
    ifnone
        (M2 => OA2) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BEM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEM8RA (M0, M1, M2, OA1, OA2, Z);
  input M0, M1, M2;
  output OA1, OA2, Z;

    and SMC_I0(OUT0, M0, M1);
    not SMC_I1(M2_bar, M2);
    buf SMC_I2(OUT1, M2_bar);
    or SMC_I3(OA1, OUT0, OUT1);

    not SMC_I4(M0_bar, M0);
    not SMC_I5(M1_bar, M1);
    and SMC_I6(OUT2, M0_bar, M1_bar);
    buf SMC_I7(OUT3, M2);
    or SMC_I8(OA2, OUT2, OUT3);

    xnor SMC_I9(Z, M0, M1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> OA1
    (M0 => OA1) = (0.0, 0.0);

    // arc M0 --> OA2
    (M0 => OA2) = (0.0, 0.0);

    // arc M0 --> Z
    if (M1===1'b0 && M2===1'b0)
        (M0 => Z) = (0.0, 0.0);
    if (M1===1'b0 && M2===1'b1)
        (M0 => Z) = (0.0, 0.0);
    if (M1===1'b1 && M2===1'b0)
        (M0 => Z) = (0.0, 0.0);
    if (M1===1'b1 && M2===1'b1)
        (M0 => Z) = (0.0, 0.0);
    ifnone
        (M0 => Z) = (0.0, 0.0);

    // arc M1 --> OA1
    (M1 => OA1) = (0.0, 0.0);

    // arc M1 --> OA2
    (M1 => OA2) = (0.0, 0.0);

    // arc M1 --> Z
    if (M0===1'b0 && M2===1'b0)
        (M1 => Z) = (0.0, 0.0);
    if (M0===1'b0 && M2===1'b1)
        (M1 => Z) = (0.0, 0.0);
    if (M0===1'b1 && M2===1'b0)
        (M1 => Z) = (0.0, 0.0);
    if (M0===1'b1 && M2===1'b1)
        (M1 => Z) = (0.0, 0.0);
    ifnone
        (M1 => Z) = (0.0, 0.0);

    // arc M2 --> OA1
    if (M0===1'b0 && M1===1'b0)
        (M2 => OA1) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1)
        (M2 => OA1) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0)
        (M2 => OA1) = (0.0, 0.0);
    ifnone
        (M2 => OA1) = (0.0, 0.0);

    // arc M2 --> OA2
    if (M0===1'b0 && M1===1'b1)
        (M2 => OA2) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0)
        (M2 => OA2) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1)
        (M2 => OA2) = (0.0, 0.0);
    ifnone
        (M2 => OA2) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BEM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEMXBM2R ( PB, M0, M1, OA1, OA2, Z );
   input M0, M1, OA1, OA2, Z;
   output PB;
      BEMXB_UDP5(PB, M0, M1, OA1, OA2, Z);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> PB
    if (M1===1'b0 && OA1===1'b0 && OA2===1'b1 && Z===1'b1)
        (M0 => PB) = (0.0, 0.0);
    if (M1===1'b0 && OA1===1'b1 && OA2===1'b0 && Z===1'b1)
        (M0 => PB) = (0.0, 0.0);
    if (M1===1'b1 && OA1===1'b0 && OA2===1'b1 && Z===1'b1)
        (M0 => PB) = (0.0, 0.0);
    if (M1===1'b1 && OA1===1'b1 && OA2===1'b0 && Z===1'b1)
        (M0 => PB) = (0.0, 0.0);
    ifnone
        (M0 => PB) = (0.0, 0.0);

    // arc M1 --> PB
    if (M0===1'b0 && OA1===1'b0 && OA2===1'b1 && Z===1'b0)
        (M1 => PB) = (0.0, 0.0);
    if (M0===1'b0 && OA1===1'b1 && OA2===1'b0 && Z===1'b0)
        (M1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && OA1===1'b0 && OA2===1'b1 && Z===1'b0)
        (M1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && OA1===1'b1 && OA2===1'b0 && Z===1'b0)
        (M1 => PB) = (0.0, 0.0);
    ifnone
        (M1 => PB) = (0.0, 0.0);

    // arc OA1 --> PB
    if (M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1)
        (OA1 => PB) = (0.0, 0.0);
    ifnone
        (OA1 => PB) = (0.0, 0.0);

    // arc OA2 --> PB
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
        (OA2 => PB) = (0.0, 0.0);
    ifnone
        (OA2 => PB) = (0.0, 0.0);

    // arc Z --> PB
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1)
        (Z => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0)
        (Z => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1)
        (Z => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0)
        (Z => PB) = (0.0, 0.0);
    ifnone
        (Z => PB) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BEMXBM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEMXBM4R ( PB, M0, M1, OA1, OA2, Z );
   input M0, M1, OA1, OA2, Z;
   output PB;
      BEMXB_UDP5(PB, M0, M1, OA1, OA2, Z);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> PB
    if (M1===1'b0 && OA1===1'b0 && OA2===1'b1 && Z===1'b1)
        (M0 => PB) = (0.0, 0.0);
    if (M1===1'b0 && OA1===1'b1 && OA2===1'b0 && Z===1'b1)
        (M0 => PB) = (0.0, 0.0);
    if (M1===1'b1 && OA1===1'b0 && OA2===1'b1 && Z===1'b1)
        (M0 => PB) = (0.0, 0.0);
    if (M1===1'b1 && OA1===1'b1 && OA2===1'b0 && Z===1'b1)
        (M0 => PB) = (0.0, 0.0);
    ifnone
        (M0 => PB) = (0.0, 0.0);

    // arc M1 --> PB
    if (M0===1'b0 && OA1===1'b0 && OA2===1'b1 && Z===1'b0)
        (M1 => PB) = (0.0, 0.0);
    if (M0===1'b0 && OA1===1'b1 && OA2===1'b0 && Z===1'b0)
        (M1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && OA1===1'b0 && OA2===1'b1 && Z===1'b0)
        (M1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && OA1===1'b1 && OA2===1'b0 && Z===1'b0)
        (M1 => PB) = (0.0, 0.0);
    ifnone
        (M1 => PB) = (0.0, 0.0);

    // arc OA1 --> PB
    if (M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
        (OA1 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1)
        (OA1 => PB) = (0.0, 0.0);
    ifnone
        (OA1 => PB) = (0.0, 0.0);

    // arc OA2 --> PB
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
        (OA2 => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
        (OA2 => PB) = (0.0, 0.0);
    ifnone
        (OA2 => PB) = (0.0, 0.0);

    // arc Z --> PB
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1)
        (Z => PB) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0)
        (Z => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1)
        (Z => PB) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0)
        (Z => PB) = (0.0, 0.0);
    ifnone
        (Z => PB) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BEMXBM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEMXM2RA ( P, M0, M1, OA1, OA2, Z );
   input M0, M1, OA1, OA2, Z;
   output P;
      BEMX_UDP5(P, M0, M1, OA1, OA2, Z);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> P
    if (M1===1'b0 && OA1===1'b0 && OA2===1'b1 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    if (M1===1'b0 && OA1===1'b1 && OA2===1'b0 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    if (M1===1'b1 && OA1===1'b0 && OA2===1'b1 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    if (M1===1'b1 && OA1===1'b1 && OA2===1'b0 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    ifnone
        (M0 => P) = (0.0, 0.0);

    // arc M1 --> P
    if (M0===1'b0 && OA1===1'b0 && OA2===1'b1 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    if (M0===1'b0 && OA1===1'b1 && OA2===1'b0 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    if (M0===1'b1 && OA1===1'b0 && OA2===1'b1 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    if (M0===1'b1 && OA1===1'b1 && OA2===1'b0 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    ifnone
        (M1 => P) = (0.0, 0.0);

    // arc OA1 --> P
    if (M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    ifnone
        (OA1 => P) = (0.0, 0.0);

    // arc OA2 --> P
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    ifnone
        (OA2 => P) = (0.0, 0.0);

    // arc Z --> P
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1)
        (Z => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0)
        (Z => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1)
        (Z => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0)
        (Z => P) = (0.0, 0.0);
    ifnone
        (Z => P) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BEMXM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEMXM4RA ( P, M0, M1, OA1, OA2, Z );
   input M0, M1, OA1, OA2, Z;
   output P;
      BEMX_UDP5(P, M0, M1, OA1, OA2, Z);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> P
    if (M1===1'b0 && OA1===1'b0 && OA2===1'b1 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    if (M1===1'b0 && OA1===1'b1 && OA2===1'b0 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    if (M1===1'b1 && OA1===1'b0 && OA2===1'b1 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    if (M1===1'b1 && OA1===1'b1 && OA2===1'b0 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    ifnone
        (M0 => P) = (0.0, 0.0);

    // arc M1 --> P
    if (M0===1'b0 && OA1===1'b0 && OA2===1'b1 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    if (M0===1'b0 && OA1===1'b1 && OA2===1'b0 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    if (M0===1'b1 && OA1===1'b0 && OA2===1'b1 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    if (M0===1'b1 && OA1===1'b1 && OA2===1'b0 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    ifnone
        (M1 => P) = (0.0, 0.0);

    // arc OA1 --> P
    if (M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    ifnone
        (OA1 => P) = (0.0, 0.0);

    // arc OA2 --> P
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    ifnone
        (OA2 => P) = (0.0, 0.0);

    // arc Z --> P
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1)
        (Z => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0)
        (Z => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1)
        (Z => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0)
        (Z => P) = (0.0, 0.0);
    ifnone
        (Z => P) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BEMXM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BEMXM8RA ( P, M0, M1, OA1, OA2, Z );
   input M0, M1, OA1, OA2, Z;
   output P;
      BEMX_UDP5(P, M0, M1, OA1, OA2, Z);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc M0 --> P
    if (M1===1'b0 && OA1===1'b0 && OA2===1'b1 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    if (M1===1'b0 && OA1===1'b1 && OA2===1'b0 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    if (M1===1'b1 && OA1===1'b0 && OA2===1'b1 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    if (M1===1'b1 && OA1===1'b1 && OA2===1'b0 && Z===1'b1)
        (M0 => P) = (0.0, 0.0);
    ifnone
        (M0 => P) = (0.0, 0.0);

    // arc M1 --> P
    if (M0===1'b0 && OA1===1'b0 && OA2===1'b1 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    if (M0===1'b0 && OA1===1'b1 && OA2===1'b0 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    if (M0===1'b1 && OA1===1'b0 && OA2===1'b1 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    if (M0===1'b1 && OA1===1'b1 && OA2===1'b0 && Z===1'b0)
        (M1 => P) = (0.0, 0.0);
    ifnone
        (M1 => P) = (0.0, 0.0);

    // arc OA1 --> P
    if (M0===1'b0 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b0 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA2===1'b1 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b0 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b0)
        (OA1 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b1 && OA2===1'b1 && Z===1'b1)
        (OA1 => P) = (0.0, 0.0);
    ifnone
        (OA1 => P) = (0.0, 0.0);

    // arc OA2 --> P
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b0 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b0 && OA1===1'b1 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && Z===1'b1)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && Z===1'b0)
        (OA2 => P) = (0.0, 0.0);
    ifnone
        (OA2 => P) = (0.0, 0.0);

    // arc Z --> P
    if (M0===1'b0 && M1===1'b1 && OA1===1'b0 && OA2===1'b1)
        (Z => P) = (0.0, 0.0);
    if (M0===1'b0 && M1===1'b1 && OA1===1'b1 && OA2===1'b0)
        (Z => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b0 && OA2===1'b1)
        (Z => P) = (0.0, 0.0);
    if (M0===1'b1 && M1===1'b0 && OA1===1'b1 && OA2===1'b0)
        (Z => P) = (0.0, 0.0);
    ifnone
        (Z => P) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BEMXM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BHDM1R (Z);
  inout Z;

    // Busholder.
  wire io_wire;

  buf(weak0,weak1) SMC_I0(Z, io_wire);
  buf              SMC_I1(io_wire, Z);

  `ifdef functional // functional //

  `else // functional //

  specify




  endspecify

  `endif // functional //
endmodule     // BHDM1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM10R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM10R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM12R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM14R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM14R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM16R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM16R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM18R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM18R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM20R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM20R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM22RA (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM22RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM24R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM24R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM26RA (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM26RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM2R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM32RA (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM32RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM3R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM40RA (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM40RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM48RA (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM48RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM4R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM5R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM5R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM6R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFM8R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // BUFM8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM0R (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM12R (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM16R (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM16R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM1R (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM20R (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM20R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM22RA (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM22RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM24RA (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM24RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM2R (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM32RA (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM32RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM3R (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM40RA (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM40RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM48RA (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM48RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM4R (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM6R (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module BUFTM8R (A, E, Z);
  input A, E;
  output Z;

    buf SMC_I0(SMC_DIN0, A);

    not SMC_I1(SMC_ZEN0, E);


    bufif0 SMC_I2(Z, SMC_DIN0, SMC_ZEN0);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0,
        0.0,
        0.0,
        0.0,
        0.0,
        0.0);



  endspecify

  `endif // functional //
endmodule     // BUFTM8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M12R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M16RA (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M2R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M3R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M4R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M6R (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKAN2M8RA (A, B, Z);
  input A, B;
  output Z;

    and SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKAN2M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM12R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM16R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM16R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM1R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM20R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM20R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM22RA (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM22RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM24R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM24R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM26RA (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM26RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM2R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM32R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM32R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM3R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM40R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM40R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM48R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM48R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM4R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM6R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKBUFM8R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKBUFM8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM12R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM16R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM16R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM1R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM20R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM20R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM22RA (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM22RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM24R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM24R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM26RA (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM26RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM2R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM32R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM32R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM3R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM40R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM40R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM48R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM48R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM4R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM6R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKINVM8R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKINVM8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M12R (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M16RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M2R (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M3R (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M4R (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M6R (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKMUX2M8R (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKMUX2M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKND2M12R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKND2M12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKND2M16RA (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKND2M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKND2M2R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKND2M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKND2M4R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKND2M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKND2M6RA (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKND2M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKND2M8R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKND2M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKXOR2M12RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKXOR2M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKXOR2M1RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKXOR2M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKXOR2M2RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKXOR2M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKXOR2M4RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKXOR2M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module CKXOR2M8RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // CKXOR2M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL1M1R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // DEL1M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL1M4R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // DEL1M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL2M1R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // DEL2M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL2M4R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // DEL2M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL3M1R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // DEL3M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL3M4R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // DEL3M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL4M1R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // DEL4M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DEL4M4R (A, Z);
  input A;
  output Z;

    buf SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // DEL4M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFAQM1RA (A, B, CK, Q);
  input A, B, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(SMC_NS_IN, A, B);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: B )) = (0.0, 0.0);



    // setup
    $setup( posedge A, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge B, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge A, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge B, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge A, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge B, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge A, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge B, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFAQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFAQM2RA (A, B, CK, Q);
  input A, B, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(SMC_NS_IN, A, B);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: B )) = (0.0, 0.0);



    // setup
    $setup( posedge A, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge B, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge A, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge B, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge A, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge B, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge A, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge B, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFAQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFAQM4RA (A, B, CK, Q);
  input A, B, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(SMC_NS_IN, A, B);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: B )) = (0.0, 0.0);



    // setup
    $setup( posedge A, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge B, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge A, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge B, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge A, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge B, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge A, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge B, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFAQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFAQM6RA (A, B, CK, Q);
  input A, B, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(SMC_NS_IN, A, B);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: B )) = (0.0, 0.0);



    // setup
    $setup( posedge A, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge B, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge A, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge B, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge A, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge B, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge A, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge B, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFAQM6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFAQM8RA (A, B, CK, Q);
  input A, B, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(SMC_NS_IN, A, B);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: B )) = (0.0, 0.0);



    // setup
    $setup( posedge A, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge B, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge A, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge B, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge A, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge B, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge A, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge B, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFAQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCM1RA (D, CKB, Q, QB);
  input D, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CKB-hl ()
    $setup(posedge D, negedge CKB, 0.0, notifier);

    // setup D-hl CKB-hl ()
    $setup(negedge D, negedge CKB, 0.0, notifier);

    // hold D-lh CKB-hl ()
    $hold(negedge CKB, posedge D, 0.0, notifier);

    // hold D-hl CKB-hl ()
    $hold(negedge CKB, negedge D, 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCM2RA (D, CKB, Q, QB);
  input D, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CKB-hl ()
    $setup(posedge D, negedge CKB, 0.0, notifier);

    // setup D-hl CKB-hl ()
    $setup(negedge D, negedge CKB, 0.0, notifier);

    // hold D-lh CKB-hl ()
    $hold(negedge CKB, posedge D, 0.0, notifier);

    // hold D-hl CKB-hl ()
    $hold(negedge CKB, negedge D, 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCM4RA (D, CKB, Q, QB);
  input D, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CKB-hl ()
    $setup(posedge D, negedge CKB, 0.0, notifier);

    // setup D-hl CKB-hl ()
    $setup(negedge D, negedge CKB, 0.0, notifier);

    // hold D-lh CKB-hl ()
    $hold(negedge CKB, posedge D, 0.0, notifier);

    // hold D-hl CKB-hl ()
    $hold(negedge CKB, negedge D, 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCM8RA (D, CKB, Q, QB);
  input D, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CKB-hl ()
    $setup(posedge D, negedge CKB, 0.0, notifier);

    // setup D-hl CKB-hl ()
    $setup(negedge D, negedge CKB, 0.0, notifier);

    // hold D-lh CKB-hl ()
    $hold(negedge CKB, posedge D, 0.0, notifier);

    // hold D-hl CKB-hl ()
    $hold(negedge CKB, negedge D, 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(negedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQM1RA (D, CKB, Q);
  input D, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB, 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB, 0.0, notifier );

    // hold
    $hold( negedge CKB, negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB, posedge D, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQM2RA (D, CKB, Q);
  input D, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB, 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB, 0.0, notifier );

    // hold
    $hold( negedge CKB, negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB, posedge D, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQM4RA (D, CKB, Q);
  input D, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB, 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB, 0.0, notifier );

    // hold
    $hold( negedge CKB, negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB, posedge D, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQM8RA (D, CKB, Q);
  input D, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB, 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB, 0.0, notifier );

    // hold
    $hold( negedge CKB, negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB, posedge D, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQRM1RA (D, RB, CKB, Q);
  input D, RB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKBDhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQRM2RA (D, RB, CKB, Q);
  input D, RB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKBDhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQRM4RA (D, RB, CKB, Q);
  input D, RB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKBDhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQRM8RA (D, RB, CKB, Q);
  input D, RB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKBDhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQRSM1RA (D, RB, SB, CKB, Q);
  input D, RB, SB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKBDhl, RB, SB);

    buf SMC_I4(shcheckCKBRBhl, SB);

    buf SMC_I5(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQRSM2RA (D, RB, SB, CKB, Q);
  input D, RB, SB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKBDhl, RB, SB);

    buf SMC_I4(shcheckCKBRBhl, SB);

    buf SMC_I5(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQRSM4RA (D, RB, SB, CKB, Q);
  input D, RB, SB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKBDhl, RB, SB);

    buf SMC_I4(shcheckCKBRBhl, SB);

    buf SMC_I5(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQRSM8RA (D, RB, SB, CKB, Q);
  input D, RB, SB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKBDhl, RB, SB);

    buf SMC_I4(shcheckCKBRBhl, SB);

    buf SMC_I5(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQSM1RA (D, SB, CKB, Q);
  input D, SB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKBDhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQSM2RA (D, SB, CKB, Q);
  input D, SB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKBDhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQSM4RA (D, SB, CKB, Q);
  input D, SB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKBDhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCQSM8RA (D, SB, CKB, Q);
  input D, SB, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKBDhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCQSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCRM1RA (D, RB, CKB, Q, QB);
  input D, RB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKBDhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCRM2RA (D, RB, CKB, Q, QB);
  input D, RB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKBDhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCRM4RA (D, RB, CKB, Q, QB);
  input D, RB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKBDhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCRM8RA (D, RB, CKB, Q, QB);
  input D, RB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKBDhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCRSM1RA (D, RB, SB, CKB, Q, QB);
  input D, RB, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKBDhl, RB, SB);

    buf SMC_I6(shcheckCKBRBhl, SB);

    buf SMC_I7(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCRSM2RA (D, RB, SB, CKB, Q, QB);
  input D, RB, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKBDhl, RB, SB);

    buf SMC_I6(shcheckCKBRBhl, SB);

    buf SMC_I7(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCRSM4RA (D, RB, SB, CKB, Q, QB);
  input D, RB, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKBDhl, RB, SB);

    buf SMC_I6(shcheckCKBRBhl, SB);

    buf SMC_I7(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCRSM8RA (D, RB, SB, CKB, Q, QB);
  input D, RB, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKBDhl, RB, SB);

    buf SMC_I6(shcheckCKBRBhl, SB);

    buf SMC_I7(shcheckCKBSBhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCSM1RA (D, SB, CKB, Q, QB);
  input D, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKBDhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCSM2RA (D, SB, CKB, Q, QB);
  input D, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKBDhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCSM4RA (D, SB, CKB, Q, QB);
  input D, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKBDhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFCSM8RA (D, SB, CKB, Q, QB);
  input D, SB, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(D), .clk(SMC_CK_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKBDhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFCSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEM1RA (D, E, CK, Q, QB);
  input D, E, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEM2RA (D, E, CK, Q, QB);
  input D, E, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEM4RA (D, E, CK, Q, QB);
  input D, E, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEM8RA (D, E, CK, Q, QB);
  input D, E, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQBM1RA (D, E, CK, QB);
  input D, E, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, E);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQBM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQBM2RA (D, E, CK, QB);
  input D, E, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, E);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQBM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQBM4RA (D, E, CK, QB);
  input D, E, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, E);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQBM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQBM8RA (D, E, CK, QB);
  input D, E, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, E);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh (E)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // hold D-hl CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQBM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQM0RA (D, E, CK, Q);
  input D, E, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( posedge E, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQM0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQM1RA (D, E, CK, Q);
  input D, E, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( posedge E, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQM2RA (D, E, CK, Q);
  input D, E, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( posedge E, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQM4RA (D, E, CK, Q);
  input D, E, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( posedge E, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQM8RA (D, E, CK, Q);
  input D, E, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, E);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( posedge E, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQRM1RA (D, E, RB, CK, Q);
  input D, E, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, E, RB);

    buf SMC_I4(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQRM2RA (D, E, RB, CK, Q);
  input D, E, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, E, RB);

    buf SMC_I4(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQRM4RA (D, E, RB, CK, Q);
  input D, E, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, E, RB);

    buf SMC_I4(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQRM8RA (D, E, RB, CK, Q);
  input D, E, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, E, RB);

    buf SMC_I4(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQZRM1RA (D, E, RB, CK, Q);
  input D, E, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    DFEQZR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, E, RB);

    buf SMC_I4(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQZRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQZRM2RA (D, E, RB, CK, Q);
  input D, E, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    DFEQZR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, E, RB);

    buf SMC_I4(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQZRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQZRM4RA (D, E, RB, CK, Q);
  input D, E, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    DFEQZR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, E, RB);

    buf SMC_I4(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQZRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEQZRM8RA (D, E, RB, CK, Q);
  input D, E, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    DFEQZR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckCKDlh, E, RB);

    buf SMC_I4(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEQZRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFERM1RA (D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKDlh, E, RB);

    buf SMC_I6(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFERM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFERM2RA (D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKDlh, E, RB);

    buf SMC_I6(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFERM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFERM4RA (D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKDlh, E, RB);

    buf SMC_I6(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFERM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFERM8RA (D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D, SMC_IQ, E);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKDlh, E, RB);

    buf SMC_I6(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFERM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEZRM1RA (D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    DFEZR_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKDlh, E, RB);

    buf SMC_I6(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && E===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && E===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (RB)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (RB)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 0.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 0.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEZRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEZRM2RA (D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    DFEZR_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKDlh, E, RB);

    buf SMC_I6(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && E===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && E===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (RB)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (RB)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 0.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 0.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEZRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEZRM4RA (D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    DFEZR_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKDlh, E, RB);

    buf SMC_I6(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && E===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && E===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (RB)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (RB)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 0.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 0.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEZRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFEZRM8RA (D, E, RB, CK, Q, QB);
  input D, E, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    DFEZR_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckCKDlh, E, RB);

    buf SMC_I6(shcheckCKElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && E===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && E===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (RB)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (RB)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 0.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 0.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFEZRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFM1RA (D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFM2RA (D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFM4RA (D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFM8RA (D, CK, Q, QB);
  input D, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFMM1RA (D1, D2, S, CK, Q, QB);
  input D1, D2, S, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D1, D2, S);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKD1lh, S);

    not SMC_I6(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFMM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFMM2RA (D1, D2, S, CK, Q, QB);
  input D1, D2, S, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D1, D2, S);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKD1lh, S);

    not SMC_I6(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFMM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFMM4RA (D1, D2, S, CK, Q, QB);
  input D1, D2, S, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D1, D2, S);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKD1lh, S);

    not SMC_I6(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFMM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFMM8RA (D1, D2, S, CK, Q, QB);
  input D1, D2, S, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, D1, D2, S);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckCKD1lh, S);

    not SMC_I6(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFMM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFMQM1RA (D1, D2, S, CK, Q);
  input D1, D2, S, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D1, D2, S);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKD1lh, S);

    not SMC_I4(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFMQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFMQM2RA (D1, D2, S, CK, Q);
  input D1, D2, S, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D1, D2, S);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKD1lh, S);

    not SMC_I4(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFMQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFMQM4RA (D1, D2, S, CK, Q);
  input D1, D2, S, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D1, D2, S);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKD1lh, S);

    not SMC_I4(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFMQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFMQM8RA (D1, D2, S, CK, Q);
  input D1, D2, S, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, D1, D2, S);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKD1lh, S);

    not SMC_I4(shcheckCKD2lh, S);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFMQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBM1RA (D, CK, QB);
  input D, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBM2RA (D, CK, QB);
  input D, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBM4RA (D, CK, QB);
  input D, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBM8RA (D, CK, QB);
  input D, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBRM1RA (D, RB, CK, QB);
  input D, RB, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBRM2RA (D, RB, CK, QB);
  input D, RB, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBRM4RA (D, RB, CK, QB);
  input D, RB, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQBRM8RA (D, RB, CK, QB);
  input D, RB, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckCKDlh, RB);


  specify


    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQBRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQM1RA (D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQM2RA (D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQM4RA (D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQM8RA (D, CK, Q);
  input D, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRM1RA (D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I2(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRM2RA (D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I2(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRM4RA (D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I2(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRM8RA (D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I2(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRSM1RA (D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB)
          );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I2(shcheckCKDlh, RB, SB);

    buf SMC_I3(shcheckCKRBlh, SB);

    buf SMC_I4(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRSM2RA (D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB)
          );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I2(shcheckCKDlh, RB, SB);

    buf SMC_I3(shcheckCKRBlh, SB);

    buf SMC_I4(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRSM4RA (D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB)
          );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I2(shcheckCKDlh, RB, SB);

    buf SMC_I3(shcheckCKRBlh, SB);

    buf SMC_I4(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQRSM8RA (D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB)
          );

  `else // functional //

    dff_p0 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I2(shcheckCKDlh, RB, SB);

    buf SMC_I3(shcheckCKRBlh, SB);

    buf SMC_I4(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQSM1RA (D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I2(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQSM2RA (D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I2(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQSM4RA (D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I2(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQSM8RA (D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;


  `ifdef functional // functional //

    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I0(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I1(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I2(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZRM1RA (D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(SMC_NS_IN, D, RB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZRM2RA (D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(SMC_NS_IN, D, RB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZRM4RA (D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(SMC_NS_IN, D, RB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZRM8RA (D, RB, CK, Q);
  input D, RB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(SMC_NS_IN, D, RB);


  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZRSM1RA (D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SB_bar, SB);
    and SMC_I1(OUT0, RB, SB_bar);
    and SMC_I2(OUT1, D, RB);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(shcheckCKDlh, RB);

    buf SMC_I7(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZRSM2RA (D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SB_bar, SB);
    and SMC_I1(OUT0, RB, SB_bar);
    and SMC_I2(OUT1, D, RB);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(shcheckCKDlh, RB);

    buf SMC_I7(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZRSM4RA (D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SB_bar, SB);
    and SMC_I1(OUT0, RB, SB_bar);
    and SMC_I2(OUT1, D, RB);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(shcheckCKDlh, RB);

    buf SMC_I7(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZRSM8RA (D, RB, SB, CK, Q);
  input D, RB, SB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SB_bar, SB);
    and SMC_I1(OUT0, RB, SB_bar);
    and SMC_I2(OUT1, D, RB);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I6(shcheckCKDlh, RB);

    buf SMC_I7(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZSM1RA (D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(D_bar, D);
    nand SMC_I1(SMC_NS_IN, D_bar, SB);


  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZSM2RA (D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(D_bar, D);
    nand SMC_I1(SMC_NS_IN, D_bar, SB);


  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZSM4RA (D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(D_bar, D);
    nand SMC_I1(SMC_NS_IN, D_bar, SB);


  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFQZSM8RA (D, SB, CK, Q);
  input D, SB, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(D_bar, D);
    nand SMC_I1(SMC_NS_IN, D_bar, SB);


  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFQZSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRM1RA (D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRM2RA (D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRM4RA (D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRM8RA (D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(1'b1),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (RB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (RB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRSM1RA (D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckCKDlh, RB, SB);

    buf SMC_I5(shcheckCKRBlh, SB);

    buf SMC_I6(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRSM2RA (D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckCKDlh, RB, SB);

    buf SMC_I5(shcheckCKRBlh, SB);

    buf SMC_I6(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRSM4RA (D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckCKDlh, RB, SB);

    buf SMC_I5(shcheckCKRBlh, SB);

    buf SMC_I6(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFRSM8RA (D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB)
          );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(RB), .preset(SB),
          .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckCKDlh, RB, SB);

    buf SMC_I5(shcheckCKRBlh, SB);

    buf SMC_I6(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFSM1RA (D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFSM2RA (D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFSM4RA (D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFSM8RA (D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(D), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckCKDlh, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (CK===1'b0 && D===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh CK-lh (SB)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (SB)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRM1RA (D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(SMC_NS_IN, D, RB);


  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    if (D===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 0.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 0.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRM2RA (D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(SMC_NS_IN, D, RB);


  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    if (D===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 0.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 0.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRM4RA (D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(SMC_NS_IN, D, RB);


  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    if (D===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 0.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 0.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRM8RA (D, RB, CK, Q, QB);
  input D, RB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(SMC_NS_IN, D, RB);


  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    if (D===1'b0 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh ()
    $setup(negedge D, posedge CK, 0.0, notifier);

    // setup D-lh CK-lh ()
    $setup(posedge D, posedge CK, 0.0, notifier);

    // setup RB-hl CK-lh ()
    $setup(negedge RB, posedge CK, 0.0, notifier);

    // setup RB-lh CK-lh ()
    $setup(posedge RB, posedge CK, 0.0, notifier);

    // hold D-hl CK-lh ()
    $hold(posedge CK, negedge D, 0.0, notifier);

    // hold D-lh CK-lh ()
    $hold(posedge CK, posedge D, 0.0, notifier);

    // hold RB-hl CK-lh ()
    $hold(posedge CK, negedge RB, 0.0, notifier);

    // hold RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRSM1RA (D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(SB_bar, SB);
    and SMC_I2(OUT0, RB, SB_bar);
    and SMC_I3(OUT1, D, RB);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I8(shcheckCKDlh, RB);

    buf SMC_I9(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRSM2RA (D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(SB_bar, SB);
    and SMC_I2(OUT0, RB, SB_bar);
    and SMC_I3(OUT1, D, RB);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I8(shcheckCKDlh, RB);

    buf SMC_I9(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRSM4RA (D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(SB_bar, SB);
    and SMC_I2(OUT0, RB, SB_bar);
    and SMC_I3(OUT1, D, RB);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I8(shcheckCKDlh, RB);

    buf SMC_I9(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZRSM8RA (D, RB, SB, CK, Q, QB);
  input D, RB, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(SB_bar, SB);
    and SMC_I2(OUT0, RB, SB_bar);
    and SMC_I3(OUT1, D, RB);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I8(shcheckCKDlh, RB);

    buf SMC_I9(shcheckCKSBlh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZSM1RA (D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(D_bar, D);
    nand SMC_I2(SMC_NS_IN, D_bar, SB);


  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZSM2RA (D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(D_bar, D);
    nand SMC_I2(SMC_NS_IN, D_bar, SB);


  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZSM4RA (D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(D_bar, D);
    nand SMC_I2(SMC_NS_IN, D_bar, SB);


  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module DFZSM8RA (D, SB, CK, Q, QB);
  input D, SB, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(D_bar, D);
    nand SMC_I2(SMC_NS_IN, D_bar, SB);


  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge D, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // DFZSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM0R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM10R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM10R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM12R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM14R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM14R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM16R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM16R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM18R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM18R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM1R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM20R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM20R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM22RA (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM22RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM24R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM24R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM26RA (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM26RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM2R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM32R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM32R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM3R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM40R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM40R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM48R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM48R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM4R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM5R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM5R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM6R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module INVM8R (A, Z);
  input A;
  output Z;

    not SMC_I0(Z, A);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // INVM8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACM1RA (D, GB, Q, QB);
  input D, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl GB-lh ()
    $setup(negedge D, posedge GB, 0.0, notifier);

    // setup D-lh GB-lh ()
    $setup(posedge D, posedge GB, 0.0, notifier);

    // hold D-hl GB-lh ()
    $hold(posedge GB, negedge D, 0.0, notifier);

    // hold D-lh GB-lh ()
    $hold(posedge GB, posedge D, 0.0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 0.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 0.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACM2RA (D, GB, Q, QB);
  input D, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl GB-lh ()
    $setup(negedge D, posedge GB, 0.0, notifier);

    // setup D-lh GB-lh ()
    $setup(posedge D, posedge GB, 0.0, notifier);

    // hold D-hl GB-lh ()
    $hold(posedge GB, negedge D, 0.0, notifier);

    // hold D-lh GB-lh ()
    $hold(posedge GB, posedge D, 0.0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 0.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 0.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACM4RA (D, GB, Q, QB);
  input D, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl GB-lh ()
    $setup(negedge D, posedge GB, 0.0, notifier);

    // setup D-lh GB-lh ()
    $setup(posedge D, posedge GB, 0.0, notifier);

    // hold D-hl GB-lh ()
    $hold(posedge GB, negedge D, 0.0, notifier);

    // hold D-lh GB-lh ()
    $hold(posedge GB, posedge D, 0.0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 0.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 0.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACM8RA (D, GB, Q, QB);
  input D, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl GB-lh ()
    $setup(negedge D, posedge GB, 0.0, notifier);

    // setup D-lh GB-lh ()
    $setup(posedge D, posedge GB, 0.0, notifier);

    // hold D-hl GB-lh ()
    $hold(posedge GB, negedge D, 0.0, notifier);

    // hold D-lh GB-lh ()
    $hold(posedge GB, posedge D, 0.0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 0.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 0.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQM1RA (D, GB, Q);
  input D, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB, 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB, 0.0, notifier );

    // hold
    $hold( posedge GB, negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB, posedge D, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQM2RA (D, GB, Q);
  input D, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB, 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB, 0.0, notifier );

    // hold
    $hold( posedge GB, negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB, posedge D, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQM4RA (D, GB, Q);
  input D, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB, 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB, 0.0, notifier );

    // hold
    $hold( posedge GB, negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB, posedge D, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQM8RA (D, GB, Q);
  input D, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB, 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB, 0.0, notifier );

    // hold
    $hold( posedge GB, negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB, posedge D, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQRM1RA (D, RB, GB, Q);
  input D, RB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGBDlh, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQRM2RA (D, RB, GB, Q);
  input D, RB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGBDlh, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQRM4RA (D, RB, GB, Q);
  input D, RB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGBDlh, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQRM8RA (D, RB, GB, Q);
  input D, RB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGBDlh, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQRSM1RA (D, RB, SB, GB, Q);
  input D, RB, SB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckGBDlh, RB, SB);

    buf SMC_I5(shcheckGBRBlh, SB);

    buf SMC_I6(shcheckGBSBlh, RB);

    buf SMC_I7(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB &&&
        (shcheckGBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB &&&
        (shcheckRBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB &&&
        (shcheckGBRBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge GB &&&
        (shcheckGBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge RB &&&
        (shcheckRBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge GB &&&
        (shcheckGBRBlh === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQRSM2RA (D, RB, SB, GB, Q);
  input D, RB, SB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckGBDlh, RB, SB);

    buf SMC_I5(shcheckGBRBlh, SB);

    buf SMC_I6(shcheckGBSBlh, RB);

    buf SMC_I7(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB &&&
        (shcheckGBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB &&&
        (shcheckRBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB &&&
        (shcheckGBRBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge GB &&&
        (shcheckGBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge RB &&&
        (shcheckRBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge GB &&&
        (shcheckGBRBlh === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQRSM4RA (D, RB, SB, GB, Q);
  input D, RB, SB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckGBDlh, RB, SB);

    buf SMC_I5(shcheckGBRBlh, SB);

    buf SMC_I6(shcheckGBSBlh, RB);

    buf SMC_I7(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB &&&
        (shcheckGBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB &&&
        (shcheckRBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB &&&
        (shcheckGBRBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge GB &&&
        (shcheckGBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge RB &&&
        (shcheckRBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge GB &&&
        (shcheckGBRBlh === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQRSM8RA (D, RB, SB, GB, Q);
  input D, RB, SB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckGBDlh, RB, SB);

    buf SMC_I5(shcheckGBRBlh, SB);

    buf SMC_I6(shcheckGBSBlh, RB);

    buf SMC_I7(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB &&&
        (shcheckGBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB &&&
        (shcheckRBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB &&&
        (shcheckGBRBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge GB &&&
        (shcheckGBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge RB &&&
        (shcheckRBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge GB &&&
        (shcheckGBRBlh === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQSM1RA (D, SB, GB, Q);
  input D, SB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGBDlh, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQSM2RA (D, SB, GB, Q);
  input D, SB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGBDlh, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQSM4RA (D, SB, GB, Q);
  input D, SB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGBDlh, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACQSM8RA (D, SB, GB, Q);
  input D, SB, GB;
  output Q;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGBDlh, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACQSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRM1RA (D, RB, GB, Q, QB);
  input D, RB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckGBDlh, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRM2RA (D, RB, GB, Q, QB);
  input D, RB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckGBDlh, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRM4RA (D, RB, GB, Q, QB);
  input D, RB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckGBDlh, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRM8RA (D, RB, GB, Q, QB);
  input D, RB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckGBDlh, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRSM1RA (D, RB, SB, GB, Q, QB);
  input D, RB, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckGBDlh, RB, SB);

    buf SMC_I6(shcheckGBRBlh, SB);

    buf SMC_I7(shcheckGBSBlh, RB);

    buf SMC_I8(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (D===1'b0 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (D===1'b0 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (D===1'b0 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (D===1'b0 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh GB-lh (RB&SB)
    $setup(posedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // setup D-hl GB-lh (RB&SB)
    $setup(negedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // setup SB-lh RB-lh (GB)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // hold D-lh GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        posedge D &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // hold D-hl GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        negedge D &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // hold SB-lh RB-lh (GB)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // recovery SB-lh RB-lh (GB)
    $recovery(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // recovery RB-lh GB-lh (SB)
    $recovery(posedge RB &&& (shcheckGBRBlh === 1'b1),
        posedge GB &&& (shcheckGBRBlh === 1'b1), 0.0, notifier);

    // recovery SB-lh GB-lh (RB)
    $recovery(posedge SB &&& (shcheckGBSBlh === 1'b1),
        posedge GB &&& (shcheckGBSBlh === 1'b1), 0.0, notifier);

    // removal RB-lh GB-lh (SB)
    $hold(posedge GB &&& (shcheckGBRBlh === 1'b1),
        posedge RB &&& (shcheckGBRBlh === 1'b1), 0.0, notifier);

    // removal SB-lh GB-lh (RB)
    $hold(posedge GB &&& (shcheckGBSBlh === 1'b1),
        posedge SB &&& (shcheckGBSBlh === 1'b1), 0.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 0.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 0.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRSM2RA (D, RB, SB, GB, Q, QB);
  input D, RB, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckGBDlh, RB, SB);

    buf SMC_I6(shcheckGBRBlh, SB);

    buf SMC_I7(shcheckGBSBlh, RB);

    buf SMC_I8(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (D===1'b0 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (D===1'b0 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (D===1'b0 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (D===1'b0 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh GB-lh (RB&SB)
    $setup(posedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // setup D-hl GB-lh (RB&SB)
    $setup(negedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // setup SB-lh RB-lh (GB)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // hold D-lh GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        posedge D &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // hold D-hl GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        negedge D &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // hold SB-lh RB-lh (GB)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // recovery SB-lh RB-lh (GB)
    $recovery(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // recovery RB-lh GB-lh (SB)
    $recovery(posedge RB &&& (shcheckGBRBlh === 1'b1),
        posedge GB &&& (shcheckGBRBlh === 1'b1), 0.0, notifier);

    // recovery SB-lh GB-lh (RB)
    $recovery(posedge SB &&& (shcheckGBSBlh === 1'b1),
        posedge GB &&& (shcheckGBSBlh === 1'b1), 0.0, notifier);

    // removal RB-lh GB-lh (SB)
    $hold(posedge GB &&& (shcheckGBRBlh === 1'b1),
        posedge RB &&& (shcheckGBRBlh === 1'b1), 0.0, notifier);

    // removal SB-lh GB-lh (RB)
    $hold(posedge GB &&& (shcheckGBSBlh === 1'b1),
        posedge SB &&& (shcheckGBSBlh === 1'b1), 0.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 0.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 0.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRSM4RA (D, RB, SB, GB, Q, QB);
  input D, RB, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckGBDlh, RB, SB);

    buf SMC_I6(shcheckGBRBlh, SB);

    buf SMC_I7(shcheckGBSBlh, RB);

    buf SMC_I8(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (D===1'b0 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (D===1'b0 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (D===1'b0 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (D===1'b0 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh GB-lh (RB&SB)
    $setup(posedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // setup D-hl GB-lh (RB&SB)
    $setup(negedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // setup SB-lh RB-lh (GB)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // hold D-lh GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        posedge D &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // hold D-hl GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        negedge D &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // hold SB-lh RB-lh (GB)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // recovery SB-lh RB-lh (GB)
    $recovery(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // recovery RB-lh GB-lh (SB)
    $recovery(posedge RB &&& (shcheckGBRBlh === 1'b1),
        posedge GB &&& (shcheckGBRBlh === 1'b1), 0.0, notifier);

    // recovery SB-lh GB-lh (RB)
    $recovery(posedge SB &&& (shcheckGBSBlh === 1'b1),
        posedge GB &&& (shcheckGBSBlh === 1'b1), 0.0, notifier);

    // removal RB-lh GB-lh (SB)
    $hold(posedge GB &&& (shcheckGBRBlh === 1'b1),
        posedge RB &&& (shcheckGBRBlh === 1'b1), 0.0, notifier);

    // removal SB-lh GB-lh (RB)
    $hold(posedge GB &&& (shcheckGBSBlh === 1'b1),
        posedge SB &&& (shcheckGBSBlh === 1'b1), 0.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 0.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 0.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACRSM8RA (D, RB, SB, GB, Q, QB);
  input D, RB, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I5(shcheckGBDlh, RB, SB);

    buf SMC_I6(shcheckGBRBlh, SB);

    buf SMC_I7(shcheckGBSBlh, RB);

    buf SMC_I8(shcheckRBSBlh, GB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (D===1'b0 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (D===1'b0 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (D===1'b0 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (D===1'b0 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && GB===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh GB-lh (RB&SB)
    $setup(posedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // setup D-hl GB-lh (RB&SB)
    $setup(negedge D &&& (shcheckGBDlh === 1'b1),
        posedge GB &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // setup SB-lh RB-lh (GB)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // hold D-lh GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        posedge D &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // hold D-hl GB-lh (RB&SB)
    $hold(posedge GB &&& (shcheckGBDlh === 1'b1),
        negedge D &&& (shcheckGBDlh === 1'b1), 0.0, notifier);

    // hold SB-lh RB-lh (GB)
    $hold(posedge RB &&& (shcheckRBSBlh === 1'b1),
        posedge SB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // recovery SB-lh RB-lh (GB)
    $recovery(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // recovery RB-lh GB-lh (SB)
    $recovery(posedge RB &&& (shcheckGBRBlh === 1'b1),
        posedge GB &&& (shcheckGBRBlh === 1'b1), 0.0, notifier);

    // recovery SB-lh GB-lh (RB)
    $recovery(posedge SB &&& (shcheckGBSBlh === 1'b1),
        posedge GB &&& (shcheckGBSBlh === 1'b1), 0.0, notifier);

    // removal RB-lh GB-lh (SB)
    $hold(posedge GB &&& (shcheckGBRBlh === 1'b1),
        posedge RB &&& (shcheckGBRBlh === 1'b1), 0.0, notifier);

    // removal SB-lh GB-lh (RB)
    $hold(posedge GB &&& (shcheckGBSBlh === 1'b1),
        posedge SB &&& (shcheckGBSBlh === 1'b1), 0.0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    // mpw GB-lh NS-lh ()
    $width(posedge GB, 0.0, 0, notifier);

    // mpw GB-hl NS-hl ()
    $width(negedge GB, 0.0, 0, notifier);

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACSM1RA (D, SB, GB, Q, QB);
  input D, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckGBDlh, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACSM2RA (D, SB, GB, Q, QB);
  input D, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckGBDlh, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACSM4RA (D, SB, GB, Q, QB);
  input D, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckGBDlh, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LACSM8RA (D, SB, GB, Q, QB);
  input D, SB, GB;
  output Q, QB;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, GB);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I2(.q(SMC_IQ), .d(D), .en(SMC_EN_IN), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I5(shcheckGBDlh, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc GB --> Q
    (negedge GB => ( Q +: D )) = (0.0, 0.0);

    // arc GB --> QB
    (negedge GB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge GB &&&
        (shcheckGBDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge GB &&&
        (shcheckGBDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge GB, 0.0, notifier );

    // removal
    $hold( posedge GB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge GB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge GB, 0.0, 0, notifier );

    $period( posedge GB, 0, notifier );
    $period( negedge GB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LACSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCECSM12RA (E, SE, CKB, GCK);
  input E, SE, CKB;
  output GCK;
  reg notifier;

  wire SMC_LD_IN;
    buf SMC_I0(OUT0, E);
    buf SMC_I1(OUT1, SE);
    or SMC_I2(SMC_LD_IN, OUT0, OUT1);

    not SMC_I3(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    not SMC_I6(CKB_bar, CKB);
    nand SMC_I7(GCK, CKB_bar, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> GCK
    (negedge CKB => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CKB-hl ()
    $setup(negedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup E-lh CKB-hl ()
    $setup(posedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // hold E-hl CKB-hl ()
    $hold(negedge CKB, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CKB-hl ()
    $hold(negedge CKB, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCECSM12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCECSM16RA (E, SE, CKB, GCK);
  input E, SE, CKB;
  output GCK;
  reg notifier;

  wire SMC_LD_IN;
    buf SMC_I0(OUT0, E);
    buf SMC_I1(OUT1, SE);
    or SMC_I2(SMC_LD_IN, OUT0, OUT1);

    not SMC_I3(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    not SMC_I6(CKB_bar, CKB);
    nand SMC_I7(GCK, CKB_bar, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> GCK
    (negedge CKB => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CKB-hl ()
    $setup(negedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup E-lh CKB-hl ()
    $setup(posedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // hold E-hl CKB-hl ()
    $hold(negedge CKB, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CKB-hl ()
    $hold(negedge CKB, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCECSM16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCECSM24RA (E, SE, CKB, GCK);
  input E, SE, CKB;
  output GCK;
  reg notifier;

  wire SMC_LD_IN;
    buf SMC_I0(OUT0, E);
    buf SMC_I1(OUT1, SE);
    or SMC_I2(SMC_LD_IN, OUT0, OUT1);

    not SMC_I3(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    not SMC_I6(CKB_bar, CKB);
    nand SMC_I7(GCK, CKB_bar, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> GCK
    (negedge CKB => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CKB-hl ()
    $setup(negedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup E-lh CKB-hl ()
    $setup(posedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // hold E-hl CKB-hl ()
    $hold(negedge CKB, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CKB-hl ()
    $hold(negedge CKB, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCECSM24RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCECSM2RA (E, SE, CKB, GCK);
  input E, SE, CKB;
  output GCK;
  reg notifier;

  wire SMC_LD_IN;
    buf SMC_I0(OUT0, E);
    buf SMC_I1(OUT1, SE);
    or SMC_I2(SMC_LD_IN, OUT0, OUT1);

    not SMC_I3(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    not SMC_I6(CKB_bar, CKB);
    nand SMC_I7(GCK, CKB_bar, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> GCK
    (negedge CKB => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CKB-hl ()
    $setup(negedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup E-lh CKB-hl ()
    $setup(posedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // hold E-hl CKB-hl ()
    $hold(negedge CKB, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CKB-hl ()
    $hold(negedge CKB, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCECSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCECSM32RA (E, SE, CKB, GCK);
  input E, SE, CKB;
  output GCK;
  reg notifier;

  wire SMC_LD_IN;
    buf SMC_I0(OUT0, E);
    buf SMC_I1(OUT1, SE);
    or SMC_I2(SMC_LD_IN, OUT0, OUT1);

    not SMC_I3(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    not SMC_I6(CKB_bar, CKB);
    nand SMC_I7(GCK, CKB_bar, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> GCK
    (negedge CKB => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CKB-hl ()
    $setup(negedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup E-lh CKB-hl ()
    $setup(posedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // hold E-hl CKB-hl ()
    $hold(negedge CKB, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CKB-hl ()
    $hold(negedge CKB, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCECSM32RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCECSM40RA (E, SE, CKB, GCK);
  input E, SE, CKB;
  output GCK;
  reg notifier;

  wire SMC_LD_IN;
    buf SMC_I0(OUT0, E);
    buf SMC_I1(OUT1, SE);
    or SMC_I2(SMC_LD_IN, OUT0, OUT1);

    not SMC_I3(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    not SMC_I6(CKB_bar, CKB);
    nand SMC_I7(GCK, CKB_bar, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> GCK
    (negedge CKB => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CKB-hl ()
    $setup(negedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup E-lh CKB-hl ()
    $setup(posedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // hold E-hl CKB-hl ()
    $hold(negedge CKB, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CKB-hl ()
    $hold(negedge CKB, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCECSM40RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCECSM48RA (E, SE, CKB, GCK);
  input E, SE, CKB;
  output GCK;
  reg notifier;

  wire SMC_LD_IN;
    buf SMC_I0(OUT0, E);
    buf SMC_I1(OUT1, SE);
    or SMC_I2(SMC_LD_IN, OUT0, OUT1);

    not SMC_I3(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    not SMC_I6(CKB_bar, CKB);
    nand SMC_I7(GCK, CKB_bar, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> GCK
    (negedge CKB => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CKB-hl ()
    $setup(negedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup E-lh CKB-hl ()
    $setup(posedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // hold E-hl CKB-hl ()
    $hold(negedge CKB, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CKB-hl ()
    $hold(negedge CKB, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCECSM48RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCECSM4RA (E, SE, CKB, GCK);
  input E, SE, CKB;
  output GCK;
  reg notifier;

  wire SMC_LD_IN;
    buf SMC_I0(OUT0, E);
    buf SMC_I1(OUT1, SE);
    or SMC_I2(SMC_LD_IN, OUT0, OUT1);

    not SMC_I3(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    not SMC_I6(CKB_bar, CKB);
    nand SMC_I7(GCK, CKB_bar, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> GCK
    (negedge CKB => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CKB-hl ()
    $setup(negedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup E-lh CKB-hl ()
    $setup(posedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // hold E-hl CKB-hl ()
    $hold(negedge CKB, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CKB-hl ()
    $hold(negedge CKB, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCECSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCECSM6RA (E, SE, CKB, GCK);
  input E, SE, CKB;
  output GCK;
  reg notifier;

  wire SMC_LD_IN;
    buf SMC_I0(OUT0, E);
    buf SMC_I1(OUT1, SE);
    or SMC_I2(SMC_LD_IN, OUT0, OUT1);

    not SMC_I3(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    not SMC_I6(CKB_bar, CKB);
    nand SMC_I7(GCK, CKB_bar, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> GCK
    (negedge CKB => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CKB-hl ()
    $setup(negedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup E-lh CKB-hl ()
    $setup(posedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // hold E-hl CKB-hl ()
    $hold(negedge CKB, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CKB-hl ()
    $hold(negedge CKB, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCECSM6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCECSM8RA (E, SE, CKB, GCK);
  input E, SE, CKB;
  output GCK;
  reg notifier;

  wire SMC_LD_IN;
    buf SMC_I0(OUT0, E);
    buf SMC_I1(OUT1, SE);
    or SMC_I2(SMC_LD_IN, OUT0, OUT1);

    not SMC_I3(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1));

  `else // functional //
    ldlatch_p0 SMC_I4(.q(SMC_IQ), .d(SMC_LD_IN), .en(CKB), .clear(1'b1),
        .preset(1'b1), .notifier(notifier));

  `endif // functional //

    //  output pins

    not SMC_I6(CKB_bar, CKB);
    nand SMC_I7(GCK, CKB_bar, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CKB --> GCK
    (negedge CKB => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CKB-hl ()
    $setup(negedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup E-lh CKB-hl ()
    $setup(posedge E &&&
        (SE === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-hl CKB-hl ()
    $setup(negedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-hl ()
    $setup(posedge SE &&&
        (E === 1'b0), negedge CKB, 0.0, notifier);

    // hold E-hl CKB-hl ()
    $hold(negedge CKB, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CKB-hl ()
    $hold(negedge CKB, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CKB-hl ()
    $hold(negedge CKB, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CKB-hl ()
    $hold(negedge CKB, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(posedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCECSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM12R (E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM16R (E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM16R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM20R (E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM20R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM2R (E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM3R (E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM4R (E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM6R (E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEM8R (E, CK, GCK);
  input E, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEM8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM12R (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM16R (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM16R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM20R (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM20R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM2R (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM3R (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM4R (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM6R (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPM8R (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I3(OUT0, CK, SE);
    and SMC_I4(OUT1, CK, SMC_IQ);
    or SMC_I5(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //


  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPM8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM12R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


   // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc CK --> OBS
    if (SE===1'b0)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    if (SE===1'b1)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);

    // arc E --> OBS
    if (SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM16R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


   // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc CK --> OBS
    if (SE===1'b0)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    if (SE===1'b1)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);

    // arc E --> OBS
    if (SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM16R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM20R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


   // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc CK --> OBS
    if (SE===1'b0)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    if (SE===1'b1)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);

    // arc E --> OBS
    if (SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM20R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM2R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


   // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc CK --> OBS
    if (SE===1'b0)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    if (SE===1'b1)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);

    // arc E --> OBS
    if (SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM3R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


   // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc CK --> OBS
    if (SE===1'b0)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    if (SE===1'b1)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);

    // arc E --> OBS
    if (SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM4R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


   // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc CK --> OBS
    if (SE===1'b0)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    if (SE===1'b1)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);

    // arc E --> OBS
    if (SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM6R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


   // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc CK --> OBS
    if (SE===1'b0)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    if (SE===1'b1)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);

    // arc E --> OBS
    if (SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCEPOM8R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(E), .en(SMC_EN_IN), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(OBS, SMC_IQ);

    and SMC_I4(OUT0, CK, SE);
    and SMC_I5(OUT1, CK, SMC_IQ);
    or SMC_I6(GCK, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


   // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);

    // arc CK --> OBS
    if (SE===1'b0)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    if (SE===1'b1)
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( OBS +: E )) = (0.0, 0.0);

    // arc E --> OBS
    if (SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);

    // arc SE --> GCK
    if (E===1'b0)
        (SE => GCK) = (0.0, 0.0);
    if (E===1'b1)
        (SE => GCK) = (0.0, 0.0);
    ifnone
        (SE => GCK) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E, posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E, posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E, 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E, 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCEPOM8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM12RA (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM16RA (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM24RA (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM24RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM2RA (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM32RA (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM32RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM40RA (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM40RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM48RA (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM48RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM4RA (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM6RA (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESM8RA (E, SE, CK, GCK);
  input E, SE, CK;
  output GCK;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: E )) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM12R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);

    // arc E --> OBS
    if (CK===1'b0 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b0 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM12R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM16R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);

    // arc E --> OBS
    if (CK===1'b0 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b0 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM16R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM20R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);

    // arc E --> OBS
    if (CK===1'b0 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b0 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM20R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM2R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);

    // arc E --> OBS
    if (CK===1'b0 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b0 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM3R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);

    // arc E --> OBS
    if (CK===1'b0 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b0 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM4R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);

    // arc E --> OBS
    if (CK===1'b0 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b0 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM6R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);

    // arc E --> OBS
    if (CK===1'b0 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b0 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAGCESOM8R (E, SE, CK, GCK, OBS);
  input E, SE, CK;
  output GCK, OBS;
  reg notifier;

  wire SMC_EN_IN;
    not SMC_I0(SMC_EN_IN, CK);

  wire SMC_LD_IN;
    buf SMC_I1(OUT0, E);
    buf SMC_I2(OUT1, SE);
    or SMC_I3(SMC_LD_IN, OUT0, OUT1);

    not SMC_I4(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I5(.q(SMC_IQ), .d(SMC_LD_IN), .en(SMC_EN_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    and SMC_I6(GCK, CK, SMC_IQ);

    buf SMC_I7(OBS, E);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc CK --> GCK
    if (E===1'b0 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b0 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b0)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    if (E===1'b1 && SE===1'b1)
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);
    ifnone
        (negedge CK => ( GCK +: SE )) = (0.0, 0.0);

    // arc E --> OBS
    if (CK===1'b0 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b0 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b0)
        (E => OBS) = (0.0, 0.0);
    if (CK===1'b1 && SE===1'b1)
        (E => OBS) = (0.0, 0.0);
    ifnone
        (E => OBS) = (0.0, 0.0);



    // setup E-hl CK-lh ()
    $setup(negedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup E-lh CK-lh ()
    $setup(posedge E &&&
        (SE === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE &&&
        (E === 1'b0), posedge CK, 0.0, notifier);

    // hold E-hl CK-lh ()
    $hold(posedge CK, negedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold E-lh CK-lh ()
    $hold(posedge CK, posedge E &&&
        (SE === 1'b0), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE &&&
        (E === 1'b0), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAGCESOM8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAM1RA (D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 0.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 0.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 0.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 0.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 0.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 0.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAM2RA (D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 0.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 0.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 0.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 0.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 0.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 0.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAM4RA (D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 0.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 0.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 0.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 0.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 0.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 0.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAM8RA (D, G, Q, QB);
  input D, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl G-hl ()
    $setup(negedge D, negedge G, 0.0, notifier);

    // setup D-lh G-hl ()
    $setup(posedge D, negedge G, 0.0, notifier);

    // hold D-hl G-hl ()
    $hold(negedge G, negedge D, 0.0, notifier);

    // hold D-lh G-hl ()
    $hold(negedge G, posedge D, 0.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 0.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 0.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQM1RA (D, G, Q);
  input D, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G, 0.0, notifier );

    // setup
    $setup( negedge D, negedge G, 0.0, notifier );

    // hold
    $hold( negedge G, posedge D, 0.0, notifier );

    // hold
    $hold( negedge G, negedge D, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQM2RA (D, G, Q);
  input D, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G, 0.0, notifier );

    // setup
    $setup( negedge D, negedge G, 0.0, notifier );

    // hold
    $hold( negedge G, posedge D, 0.0, notifier );

    // hold
    $hold( negedge G, negedge D, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQM4RA (D, G, Q);
  input D, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G, 0.0, notifier );

    // setup
    $setup( negedge D, negedge G, 0.0, notifier );

    // hold
    $hold( negedge G, posedge D, 0.0, notifier );

    // hold
    $hold( negedge G, negedge D, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQM8RA (D, G, Q);
  input D, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G, 0.0, notifier );

    // setup
    $setup( negedge D, negedge G, 0.0, notifier );

    // hold
    $hold( negedge G, posedge D, 0.0, notifier );

    // hold
    $hold( negedge G, negedge D, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQRM1RA (D, RB, G, Q);
  input D, RB, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckGDhl, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQRM2RA (D, RB, G, Q);
  input D, RB, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckGDhl, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQRM4RA (D, RB, G, Q);
  input D, RB, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckGDhl, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQRM8RA (D, RB, G, Q);
  input D, RB, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckGDhl, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQRSM1RA (D, RB, SB, G, Q);
  input D, RB, SB, G;
  output Q;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckGDhl, RB, SB);

    buf SMC_I4(shcheckGRBhl, SB);

    buf SMC_I5(shcheckGSBhl, RB);

    not SMC_I6(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB &&&
        (shcheckRBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G &&&
        (shcheckGRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G &&&
        (shcheckGSBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge RB &&&
        (shcheckRBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( negedge G &&&
        (shcheckGRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( negedge G &&&
        (shcheckGSBhl === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQRSM2RA (D, RB, SB, G, Q);
  input D, RB, SB, G;
  output Q;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckGDhl, RB, SB);

    buf SMC_I4(shcheckGRBhl, SB);

    buf SMC_I5(shcheckGSBhl, RB);

    not SMC_I6(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB &&&
        (shcheckRBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G &&&
        (shcheckGRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G &&&
        (shcheckGSBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge RB &&&
        (shcheckRBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( negedge G &&&
        (shcheckGRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( negedge G &&&
        (shcheckGSBhl === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQRSM4RA (D, RB, SB, G, Q);
  input D, RB, SB, G;
  output Q;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckGDhl, RB, SB);

    buf SMC_I4(shcheckGRBhl, SB);

    buf SMC_I5(shcheckGSBhl, RB);

    not SMC_I6(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB &&&
        (shcheckRBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G &&&
        (shcheckGRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G &&&
        (shcheckGSBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge RB &&&
        (shcheckRBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( negedge G &&&
        (shcheckGRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( negedge G &&&
        (shcheckGSBhl === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQRSM8RA (D, RB, SB, G, Q);
  input D, RB, SB, G;
  output Q;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I3(shcheckGDhl, RB, SB);

    buf SMC_I4(shcheckGRBhl, SB);

    buf SMC_I5(shcheckGSBhl, RB);

    not SMC_I6(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB &&&
        (shcheckRBSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G &&&
        (shcheckGRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G &&&
        (shcheckGSBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge RB &&&
        (shcheckRBSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( negedge G &&&
        (shcheckGRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( negedge G &&&
        (shcheckGSBhl === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQSM1RA (D, SB, G, Q);
  input D, SB, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckGDhl, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQSM2RA (D, SB, G, Q);
  input D, SB, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckGDhl, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQSM4RA (D, SB, G, Q);
  input D, SB, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckGDhl, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LAQSM8RA (D, SB, G, Q);
  input D, SB, G;
  output Q;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I3(shcheckGDhl, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LAQSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARM1RA (D, RB, G, Q, QB);
  input D, RB, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGDhl, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARM2RA (D, RB, G, Q, QB);
  input D, RB, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGDhl, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARM4RA (D, RB, G, Q, QB);
  input D, RB, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGDhl, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARM8RA (D, RB, G, Q, QB);
  input D, RB, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGDhl, RB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARSM1RA (D, RB, SB, G, Q, QB);
  input D, RB, SB, G;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckGDhl, RB, SB);

    buf SMC_I5(shcheckGRBhl, SB);

    buf SMC_I6(shcheckGSBhl, RB);

    not SMC_I7(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (D===1'b0 && G===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (D===1'b0 && G===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (D===1'b0 && G===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (D===1'b0 && G===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh G-hl (RB&SB)
    $setup(posedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // setup D-hl G-hl (RB&SB)
    $setup(negedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // setup SB-lh RB-lh (!G)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // hold D-lh G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        posedge D &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // hold D-hl G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        negedge D &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // hold SB-lh RB-lh (!G)
    $hold(posedge RB &&& (shcheckRBSBlh===1'b1),
        posedge SB &&& (shcheckRBSBlh===1'b1), 0.0, notifier);

    // recovery SB-lh RB-lh (!G)
    $recovery(posedge SB &&& (shcheckRBSBlh===1'b1),
        posedge RB &&& (shcheckRBSBlh===1'b1), 0.0, notifier);

    // recovery SB-lh G-hl (RB)
    $recovery(posedge SB &&& (shcheckGSBhl === 1'b1),
        negedge G &&& (shcheckGSBhl === 1'b1), 0.0, notifier);

    // recovery RB-lh G-hl (SB)
    $recovery(posedge RB &&& (shcheckGRBhl === 1'b1),
        negedge G &&& (shcheckGRBhl === 1'b1), 0.0, notifier);

    // removal SB-lh G-hl (RB)
    $hold(negedge G &&& (shcheckGSBhl === 1'b1),
        posedge SB &&& (shcheckGSBhl === 1'b1), 0.0, notifier);

    // removal RB-lh G-hl (SB)
    $hold(negedge G &&& (shcheckGRBhl === 1'b1),
        posedge RB &&& (shcheckGRBhl === 1'b1), 0.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 0.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARSM2RA (D, RB, SB, G, Q, QB);
  input D, RB, SB, G;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckGDhl, RB, SB);

    buf SMC_I5(shcheckGRBhl, SB);

    buf SMC_I6(shcheckGSBhl, RB);

    not SMC_I7(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (D===1'b0 && G===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (D===1'b0 && G===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (D===1'b0 && G===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (D===1'b0 && G===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh G-hl (RB&SB)
    $setup(posedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // setup D-hl G-hl (RB&SB)
    $setup(negedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // setup SB-lh RB-lh (!G)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // hold D-lh G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        posedge D &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // hold D-hl G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        negedge D &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // hold SB-lh RB-lh (!G)
    $hold(posedge RB &&& (shcheckRBSBlh===1'b1),
        posedge SB &&& (shcheckRBSBlh===1'b1), 0.0, notifier);

    // recovery SB-lh RB-lh (!G)
    $recovery(posedge SB &&& (shcheckRBSBlh===1'b1),
        posedge RB &&& (shcheckRBSBlh===1'b1), 0.0, notifier);

    // recovery SB-lh G-hl (RB)
    $recovery(posedge SB &&& (shcheckGSBhl === 1'b1),
        negedge G &&& (shcheckGSBhl === 1'b1), 0.0, notifier);

    // recovery RB-lh G-hl (SB)
    $recovery(posedge RB &&& (shcheckGRBhl === 1'b1),
        negedge G &&& (shcheckGRBhl === 1'b1), 0.0, notifier);

    // removal SB-lh G-hl (RB)
    $hold(negedge G &&& (shcheckGSBhl === 1'b1),
        posedge SB &&& (shcheckGSBhl === 1'b1), 0.0, notifier);

    // removal RB-lh G-hl (SB)
    $hold(negedge G &&& (shcheckGRBhl === 1'b1),
        posedge RB &&& (shcheckGRBhl === 1'b1), 0.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 0.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARSM4RA (D, RB, SB, G, Q, QB);
  input D, RB, SB, G;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckGDhl, RB, SB);

    buf SMC_I5(shcheckGRBhl, SB);

    buf SMC_I6(shcheckGSBhl, RB);

    not SMC_I7(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (D===1'b0 && G===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (D===1'b0 && G===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (D===1'b0 && G===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (D===1'b0 && G===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh G-hl (RB&SB)
    $setup(posedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // setup D-hl G-hl (RB&SB)
    $setup(negedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // setup SB-lh RB-lh (!G)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // hold D-lh G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        posedge D &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // hold D-hl G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        negedge D &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // hold SB-lh RB-lh (!G)
    $hold(posedge RB &&& (shcheckRBSBlh===1'b1),
        posedge SB &&& (shcheckRBSBlh===1'b1), 0.0, notifier);

    // recovery SB-lh RB-lh (!G)
    $recovery(posedge SB &&& (shcheckRBSBlh===1'b1),
        posedge RB &&& (shcheckRBSBlh===1'b1), 0.0, notifier);

    // recovery SB-lh G-hl (RB)
    $recovery(posedge SB &&& (shcheckGSBhl === 1'b1),
        negedge G &&& (shcheckGSBhl === 1'b1), 0.0, notifier);

    // recovery RB-lh G-hl (SB)
    $recovery(posedge RB &&& (shcheckGRBhl === 1'b1),
        negedge G &&& (shcheckGRBhl === 1'b1), 0.0, notifier);

    // removal SB-lh G-hl (RB)
    $hold(negedge G &&& (shcheckGSBhl === 1'b1),
        posedge SB &&& (shcheckGSBhl === 1'b1), 0.0, notifier);

    // removal RB-lh G-hl (SB)
    $hold(negedge G &&& (shcheckGRBhl === 1'b1),
        posedge RB &&& (shcheckGRBhl === 1'b1), 0.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 0.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LARSM8RA (D, RB, SB, G, Q, QB);
  input D, RB, SB, G;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I4(shcheckGDhl, RB, SB);

    buf SMC_I5(shcheckGRBhl, SB);

    buf SMC_I6(shcheckGSBhl, RB);

    not SMC_I7(shcheckRBSBlh, G);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (D===1'b0 && G===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && SB===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (D===1'b0 && G===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && SB===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (D===1'b0 && G===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && RB===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (D===1'b0 && G===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && G===1'b1 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b0 && RB===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && G===1'b1 && RB===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-lh G-hl (RB&SB)
    $setup(posedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // setup D-hl G-hl (RB&SB)
    $setup(negedge D &&& (shcheckGDhl === 1'b1),
        negedge G &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // setup SB-lh RB-lh (!G)
    $setup(posedge SB &&& (shcheckRBSBlh === 1'b1),
        posedge RB &&& (shcheckRBSBlh === 1'b1), 0.0, notifier);

    // hold D-lh G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        posedge D &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // hold D-hl G-hl (RB&SB)
    $hold(negedge G &&& (shcheckGDhl === 1'b1),
        negedge D &&& (shcheckGDhl === 1'b1), 0.0, notifier);

    // hold SB-lh RB-lh (!G)
    $hold(posedge RB &&& (shcheckRBSBlh===1'b1),
        posedge SB &&& (shcheckRBSBlh===1'b1), 0.0, notifier);

    // recovery SB-lh RB-lh (!G)
    $recovery(posedge SB &&& (shcheckRBSBlh===1'b1),
        posedge RB &&& (shcheckRBSBlh===1'b1), 0.0, notifier);

    // recovery SB-lh G-hl (RB)
    $recovery(posedge SB &&& (shcheckGSBhl === 1'b1),
        negedge G &&& (shcheckGSBhl === 1'b1), 0.0, notifier);

    // recovery RB-lh G-hl (SB)
    $recovery(posedge RB &&& (shcheckGRBhl === 1'b1),
        negedge G &&& (shcheckGRBhl === 1'b1), 0.0, notifier);

    // removal SB-lh G-hl (RB)
    $hold(negedge G &&& (shcheckGSBhl === 1'b1),
        posedge SB &&& (shcheckGSBhl === 1'b1), 0.0, notifier);

    // removal RB-lh G-hl (SB)
    $hold(negedge G &&& (shcheckGRBhl === 1'b1),
        posedge RB &&& (shcheckGRBhl === 1'b1), 0.0, notifier);

    // mpw G-hl NS-hl ()
    $width(negedge G, 0.0, 0, notifier);

    // mpw G-lh NS-lh ()
    $width(posedge G, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LARSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LASM1RA (D, SB, G, Q, QB);
  input D, SB, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGDhl, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LASM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LASM2RA (D, SB, G, Q, QB);
  input D, SB, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGDhl, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LASM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LASM4RA (D, SB, G, Q, QB);
  input D, SB, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGDhl, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LASM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module LASM8RA (D, SB, G, Q, QB);
  input D, SB, G;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    ldlatch_p1 SMC_I1(.q(SMC_IQ), .d(D), .en(G), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    buf SMC_I4(shcheckGDhl, SB);


  specify


    // arc D --> Q
    (D => Q) = (0.0, 0.0);

    // arc D --> QB
    (D => QB) = (0.0, 0.0);

    // arc G --> Q
    (posedge G => ( Q +: D )) = (0.0, 0.0);

    // arc G --> QB
    (posedge G => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge G &&&
        (shcheckGDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge G &&&
        (shcheckGDhl === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge G, 0.0, notifier );

    // removal
    $hold( negedge G, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge G, 0.0, 0, notifier );

    // mpw
    $width( negedge G, 0.0, 0, notifier );

    $period( posedge G, 0, notifier );
    $period( negedge G, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // LASM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAO222M1RA ( Z, A, B, C );
   input A, B, C;
   output Z;
      MAO222_UDP3(Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAO222M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAO222M2RA ( Z, A, B, C );
   input A, B, C;
   output Z;
      MAO222_UDP3(Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAO222M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAO222M4RA ( Z, A, B, C );
   input A, B, C;
   output Z;
      MAO222_UDP3(Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAO222M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAO222M8RA ( Z, A, B, C );
   input A, B, C;
   output Z;
      MAO222_UDP3(Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAO222M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI2223M1RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      MAOI2223_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI2223M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI2223M2RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      MAOI2223_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI2223M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI2223M4RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      MAOI2223_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI2223M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI2223M8RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      MAOI2223_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI2223M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI222M1RA ( Z, A, B, C );
   input A, B, C;
   output Z;
      MAOI222_UDP3(Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI222M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI222M2RA ( Z, A, B, C );
   input A, B, C;
   output Z;
      MAOI222_UDP3(Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI222M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI222M4RA ( Z, A, B, C );
   input A, B, C;
   output Z;
      MAOI222_UDP3(Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI222M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI222M8RA ( Z, A, B, C );
   input A, B, C;
   output Z;
      MAOI222_UDP3(Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI222M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI22M1RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, B1);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, B1);
    and SMC_I4(OUT2, A1_bar, B2);
    and SMC_I5(OUT3, A2_bar, B2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI22M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI22M2RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, B1);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, B1);
    and SMC_I4(OUT2, A1_bar, B2);
    and SMC_I5(OUT3, A2_bar, B2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI22M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI22M4RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, B1);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, B1);
    and SMC_I4(OUT2, A1_bar, B2);
    and SMC_I5(OUT3, A2_bar, B2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI22M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MAOI22M8RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    not SMC_I0(A1_bar, A1);
    and SMC_I1(OUT0, A1_bar, B1);
    not SMC_I2(A2_bar, A2);
    and SMC_I3(OUT1, A2_bar, B1);
    and SMC_I4(OUT2, A1_bar, B2);
    and SMC_I5(OUT3, A2_bar, B2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b1 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b1 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b1 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MAOI22M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MOAI22M1RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      MOAI22_UDP4(Z, A1, A2, B1, B2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MOAI22M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MOAI22M2RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      MOAI22_UDP4(Z, A1, A2, B1, B2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MOAI22M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MOAI22M4RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      MOAI22_UDP4(Z, A1, A2, B1, B2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MOAI22M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MOAI22M8RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;
      MOAI22_UDP4(Z, A1, A2, B1, B2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MOAI22M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M0RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M12RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M1RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M2RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M3RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M3RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M4RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M6R (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX2M8R (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(S_bar, S);
    and SMC_I1(OUT0, A, S_bar);
    and SMC_I2(OUT1, B, S);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX2M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX3M0RA ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MUX3_UDP5(Z, A, B, C, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX3M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX3M1RA ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MUX3_UDP5(Z, A, B, C, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX3M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX3M2RA ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MUX3_UDP5(Z, A, B, C, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX3M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX3M4RA ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MUX3_UDP5(Z, A, B, C, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX3M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX3M8RA ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MUX3_UDP5(Z, A, B, C, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX3M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX4M0RA ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MUX4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX4M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX4M1RA ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MUX4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX4M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX4M2RA ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MUX4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX4M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX4M4R ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MUX4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX4M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MUX4M8RA ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MUX4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MUX4M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M0RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M1RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M2RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M3RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M3RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M4RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M6RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB2M8RA (A, B, S, Z);
  input A, B, S;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(S_bar, S);
    and SMC_I2(OUT0, A_bar, S_bar);
    not SMC_I3(B_bar, B);
    and SMC_I4(OUT1, B_bar, S);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && S===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && S===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc S --> Z
    if (A===1'b0 && B===1'b1)
        (S => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (S => Z) = (0.0, 0.0);
    ifnone
        (S => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB2M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB3M0RA ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MXB3_UDP5(Z, A, B, C, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB3M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB3M1RA ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MXB3_UDP5(Z, A, B, C, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB3M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB3M2RA ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MXB3_UDP5(Z, A, B, C, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB3M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB3M4RA ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MXB3_UDP5(Z, A, B, C, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB3M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB3M8RA ( Z, A, B, C, S0, S1 );
   input A, B, C, S0, S1;
   output Z;
      MXB3_UDP5(Z, A, B, C, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && S0===1'b1 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b1 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB3M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB4M0RA ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MXB4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB4M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB4M1RA ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MXB4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB4M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB4M2RA ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MXB4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB4M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB4M4RA ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MXB4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB4M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB4M6RA ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MXB4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB4M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module MXB4M8RA ( Z, A, B, C, D, S0, S1 );
   input A, B, C, D, S0, S1;
   output Z;
      MXB4_UDP6(Z, A, B, C, D, S0, S1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b0)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1 && S0===1'b1 && S1===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1 && S0===1'b0 && S1===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && S0===1'b1 && S1===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);

    // arc S0 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S1===1'b0)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S1===1'b1)
        (S0 => Z) = (0.0, 0.0);
    ifnone
        (S0 => Z) = (0.0, 0.0);

    // arc S1 --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1 && D===1'b1 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0 && D===1'b1 && S0===1'b0)
        (S1 => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1 && D===1'b0 && S0===1'b1)
        (S1 => Z) = (0.0, 0.0);
    ifnone
        (S1 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // MXB4M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M0R (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M12RA (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M16RA (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M1R (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M2R (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M4R (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M6RA (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2B1M8R (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(NA_bar, NA);
    nand SMC_I1(Z, B, NA_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2B1M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M0R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M12RA (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M16RA (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M1R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M2R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M3R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2M3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M4R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M5R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2M5R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M6R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND2M8R (A, B, Z);
  input A, B;
  output Z;

    nand SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND2M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3B1M0R ( Z, B, C, NA );
   input B, C, NA;
   output Z;

    not (tmp1, NA);
    nand (Z, B, C, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3B1M12RA ( Z, B, C, NA );
   input B, C, NA;
   output Z;

    not (tmp1, NA);
    nand (Z, B, C, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3B1M1R ( Z, B, C, NA );
   input B, C, NA;
   output Z;

    not (tmp1, NA);
    nand (Z, B, C, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3B1M2R ( Z, B, C, NA );
   input B, C, NA;
   output Z;

    not (tmp1, NA);
    nand (Z, B, C, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3B1M4R ( Z, B, C, NA );
   input B, C, NA;
   output Z;

    not (tmp1, NA);
    nand (Z, B, C, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3B1M6RA ( Z, B, C, NA );
   input B, C, NA;
   output Z;

    not (tmp1, NA);
    nand (Z, B, C, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3B1M8RA ( Z, B, C, NA );
   input B, C, NA;
   output Z;

    not (tmp1, NA);
    nand (Z, B, C, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3B1M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3M0R ( Z, A, B, C );
   input A, B, C;
   output Z;

     nand (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3M12RA ( Z, A, B, C );
   input A, B, C;
   output Z;

     nand (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3M16RA ( Z, A, B, C );
   input A, B, C;
   output Z;

     nand (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3M1R ( Z, A, B, C );
   input A, B, C;
   output Z;

     nand (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3M2R ( Z, A, B, C );
   input A, B, C;
   output Z;

     nand (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3M3R ( Z, A, B, C );
   input A, B, C;
   output Z;

     nand (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3M3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3M4RA ( Z, A, B, C );
   input A, B, C;
   output Z;

     nand (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3M6RA ( Z, A, B, C );
   input A, B, C;
   output Z;

     nand (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND3M8RA ( Z, A, B, C );
   input A, B, C;
   output Z;

     nand (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND3M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B1M0R ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

   not (tmp1, NA);
   nand (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B1M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B1M1R ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

   not (tmp1, NA);
   nand (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B1M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B1M2R ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

   not (tmp1, NA);
   nand (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B1M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B1M4R ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

   not (tmp1, NA);
   nand (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B1M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B1M6RA ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

   not (tmp1, NA);
   nand (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B1M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B1M8RA ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

   not (tmp1, NA);
   nand (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B1M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B2M0R ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;

    not (tmp1, NA);
    not (tmp2, NB);
    nand (Z, C, D, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);

    // arc NB --> Z
    (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B2M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B2M1R ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;

    not (tmp1, NA);
    not (tmp2, NB);
    nand (Z, C, D, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);

    // arc NB --> Z
    (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B2M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B2M2R ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;

    not (tmp1, NA);
    not (tmp2, NB);
    nand (Z, C, D, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);

    // arc NB --> Z
    (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B2M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B2M4R ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;

    not (tmp1, NA);
    not (tmp2, NB);
    nand (Z, C, D, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);

    // arc NB --> Z
    (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B2M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4B2M8RA ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;

    not (tmp1, NA);
    not (tmp2, NB);
    nand (Z, C, D, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);

    // arc NB --> Z
    (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4B2M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4M0R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nand (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4M16RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nand (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4M1R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nand (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4M2R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nand (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4M4R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nand (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4M6R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nand (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module ND4M8R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nand (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // ND4M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M0R (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M12RA (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M16RA (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M1R (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M2R (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M4R (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M6RA (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2B1M8R (B, NA, Z);
  input B, NA;
  output Z;

    not SMC_I0(B_bar, B);
    and SMC_I1(Z, B_bar, NA);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2B1M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M0R (A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M12RA (A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M16RA (A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M1R (A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M2R (A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M3R (A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2M3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M4R (A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M5R (A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2M5R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M6R (A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR2M8R (A, B, Z);
  input A, B;
  output Z;

    not SMC_I0(A_bar, A);
    not SMC_I1(B_bar, B);
    and SMC_I2(Z, A_bar, B_bar);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR2M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3B1M0R ( Z, B, C, NA );
   input B, C, NA;
   output Z;

   not (tmp1, NA);
   nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3B1M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3B1M1R ( Z, B, C, NA );
   input B, C, NA;
   output Z;

   not (tmp1, NA);
   nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3B1M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3B1M2R ( Z, B, C, NA );
   input B, C, NA;
   output Z;

   not (tmp1, NA);
   nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3B1M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3B1M4R ( Z, B, C, NA );
   input B, C, NA;
   output Z;

   not (tmp1, NA);
   nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3B1M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3B1M8RA ( Z, B, C, NA );
   input B, C, NA;
   output Z;

   not (tmp1, NA);
   nor (Z, tmp1, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3B1M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3M0R ( Z, A, B, C );
   input A, B, C;
   output Z;

   nor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3M16RA ( Z, A, B, C );
   input A, B, C;
   output Z;

   nor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3M1R ( Z, A, B, C );
   input A, B, C;
   output Z;

   nor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3M2R ( Z, A, B, C );
   input A, B, C;
   output Z;

   nor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3M4R ( Z, A, B, C );
   input A, B, C;
   output Z;

   nor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3M6R ( Z, A, B, C );
   input A, B, C;
   output Z;

   nor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR3M8R ( Z, A, B, C );
   input A, B, C;
   output Z;

   nor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR3M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4B1M0R ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

  not (tmp1, NA);
  nor (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4B1M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4B1M1R ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

  not (tmp1, NA);
  nor (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4B1M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4B1M2R ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

  not (tmp1, NA);
  nor (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4B1M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4B1M4R ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

  not (tmp1, NA);
  nor (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4B1M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4B1M8RA ( Z, B, C, D, NA );
   input B, C, D, NA;
   output Z;

  not (tmp1, NA);
  nor (Z, B, C, D, tmp1);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4B1M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4B2M0R ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;

   not (tmp1, NA);
   not (tmp2, NB);
   nor (Z, C, D, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);

    // arc NB --> Z
    (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4B2M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4B2M1R ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;

   not (tmp1, NA);
   not (tmp2, NB);
   nor (Z, C, D, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);

    // arc NB --> Z
    (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4B2M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4B2M2R ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;

   not (tmp1, NA);
   not (tmp2, NB);
   nor (Z, C, D, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);

    // arc NB --> Z
    (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4B2M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4B2M4R ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;

   not (tmp1, NA);
   not (tmp2, NB);
   nor (Z, C, D, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);

    // arc NB --> Z
    (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4B2M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4B2M8RA ( Z, C, D, NA, NB );
   input C, D, NA, NB;
   output Z;

   not (tmp1, NA);
   not (tmp2, NB);
   nor (Z, C, D, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc NA --> Z
    (NA => Z) = (0.0, 0.0);

    // arc NB --> Z
    (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4B2M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4M0R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nor (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4M16RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nor (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4M1R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nor (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4M2R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nor (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4M4RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nor (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4M6R ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nor (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module NR4M8RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;

    nor (Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // NR4M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA211M12RA ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;
      OA211_UDP4(Z, A1, A2, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA211M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA211M1RA ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;
      OA211_UDP4(Z, A1, A2, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA211M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA211M2RA ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;
      OA211_UDP4(Z, A1, A2, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA211M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA211M4RA ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;
      OA211_UDP4(Z, A1, A2, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA211M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA211M6RA ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;
      OA211_UDP4(Z, A1, A2, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA211M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA211M8RA ( Z, A1, A2, B, C );
   input A1, A2, B, C;
   output Z;
      OA211_UDP4(Z, A1, A2, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA211M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M0RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA21M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M12RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA21M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M16RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA21M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M1RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA21M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M2RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA21M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M4RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA21M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M6RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA21M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA21M8RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    and SMC_I0(OUT0, A1, B);
    and SMC_I1(OUT1, A2, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA21M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA221M1RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      OA221_UDP5(Z, A1, A2, B1, B2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA221M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA221M2RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      OA221_UDP5(Z, A1, A2, B1, B2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA221M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA221M4RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      OA221_UDP5(Z, A1, A2, B1, B2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA221M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA221M8RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;
      OA221_UDP5(Z, A1, A2, B1, B2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA221M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA222M1RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      OA222_UDP6(Z, A1, A2, B1, B2, C1, C2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA222M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA222M2RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      OA222_UDP6(Z, A1, A2, B1, B2, C1, C2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA222M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA222M4RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      OA222_UDP6(Z, A1, A2, B1, B2, C1, C2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA222M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA222M8RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;
      OA222_UDP6(Z, A1, A2, B1, B2, C1, C2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA222M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M0R (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA22M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M12RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA22M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M16RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA22M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M1R (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA22M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M2R (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA22M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M4R (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA22M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M6RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA22M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA22M8RA (A1, A2, B1, B2, Z);
  input A1, A2, B1, B2;
  output Z;

    and SMC_I0(OUT0, A2, B2);
    and SMC_I1(OUT1, A1, B2);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA22M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA31M1RA (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    and SMC_I0(OUT0, A3, B);
    and SMC_I1(OUT1, A1, B);
    and SMC_I2(OUT2, A2, B);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA31M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA31M2RA (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    and SMC_I0(OUT0, A3, B);
    and SMC_I1(OUT1, A1, B);
    and SMC_I2(OUT2, A2, B);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA31M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA31M4RA (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    and SMC_I0(OUT0, A3, B);
    and SMC_I1(OUT1, A1, B);
    and SMC_I2(OUT2, A2, B);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA31M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA31M8RA (A1, A2, A3, B, Z);
  input A1, A2, A3, B;
  output Z;

    and SMC_I0(OUT0, A3, B);
    and SMC_I1(OUT1, A1, B);
    and SMC_I2(OUT2, A2, B);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA31M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA32M1RA (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    and SMC_I0(OUT0, A1, B2);
    and SMC_I1(OUT1, A3, B1);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    and SMC_I4(OUT4, A2, B2);
    and SMC_I5(OUT5, A3, B2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA32M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA32M2RA (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    and SMC_I0(OUT0, A1, B2);
    and SMC_I1(OUT1, A3, B1);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    and SMC_I4(OUT4, A2, B2);
    and SMC_I5(OUT5, A3, B2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA32M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA32M4RA (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    and SMC_I0(OUT0, A1, B2);
    and SMC_I1(OUT1, A3, B1);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    and SMC_I4(OUT4, A2, B2);
    and SMC_I5(OUT5, A3, B2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA32M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA32M8RA (A1, A2, A3, B1, B2, Z);
  input A1, A2, A3, B1, B2;
  output Z;

    and SMC_I0(OUT0, A1, B2);
    and SMC_I1(OUT1, A3, B1);
    and SMC_I2(OUT2, A1, B1);
    and SMC_I3(OUT3, A2, B1);
    and SMC_I4(OUT4, A2, B2);
    and SMC_I5(OUT5, A3, B2);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA32M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA33M1RA (A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    and SMC_I0(OUT0, A3, B1);
    and SMC_I1(OUT1, A3, B3);
    and SMC_I2(OUT2, A1, B3);
    and SMC_I3(OUT3, A1, B1);
    and SMC_I4(OUT4, A1, B2);
    and SMC_I5(OUT5, A2, B1);
    and SMC_I6(OUT6, A2, B3);
    and SMC_I7(OUT7, A2, B2);
    and SMC_I8(OUT8, A3, B2);
    or SMC_I9(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I10(OUTSUB1, OUT8);
    or SMC_I11(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA33M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA33M2RA (A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    and SMC_I0(OUT0, A3, B1);
    and SMC_I1(OUT1, A3, B3);
    and SMC_I2(OUT2, A1, B3);
    and SMC_I3(OUT3, A1, B1);
    and SMC_I4(OUT4, A1, B2);
    and SMC_I5(OUT5, A2, B1);
    and SMC_I6(OUT6, A2, B3);
    and SMC_I7(OUT7, A2, B2);
    and SMC_I8(OUT8, A3, B2);
    or SMC_I9(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I10(OUTSUB1, OUT8);
    or SMC_I11(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA33M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA33M4RA (A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    and SMC_I0(OUT0, A3, B1);
    and SMC_I1(OUT1, A3, B3);
    and SMC_I2(OUT2, A1, B3);
    and SMC_I3(OUT3, A1, B1);
    and SMC_I4(OUT4, A1, B2);
    and SMC_I5(OUT5, A2, B1);
    and SMC_I6(OUT6, A2, B3);
    and SMC_I7(OUT7, A2, B2);
    and SMC_I8(OUT8, A3, B2);
    or SMC_I9(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I10(OUTSUB1, OUT8);
    or SMC_I11(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA33M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OA33M8RA (A1, A2, A3, B1, B2, B3, Z);
  input A1, A2, A3, B1, B2, B3;
  output Z;

    and SMC_I0(OUT0, A3, B1);
    and SMC_I1(OUT1, A3, B3);
    and SMC_I2(OUT2, A1, B3);
    and SMC_I3(OUT3, A1, B1);
    and SMC_I4(OUT4, A1, B2);
    and SMC_I5(OUT5, A2, B1);
    and SMC_I6(OUT6, A2, B3);
    and SMC_I7(OUT7, A2, B2);
    and SMC_I8(OUT8, A3, B2);
    or SMC_I9(OUTSUB0, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5, OUT6, OUT7);
    or SMC_I10(OUTSUB1, OUT8);
    or SMC_I11(Z, OUTSUB0, OUTSUB1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OA33M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211B100M0R (A1, B, C, NA2, Z);
  input A1, B, C, NA2;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(B_bar, B);
    buf SMC_I3(OUT1, B_bar);
    not SMC_I4(A1_bar, A1);
    and SMC_I5(OUT2, A1_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && C===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && C===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && C===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && B===1'b1 && NA2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && B===1'b1 && NA2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && B===1'b1 && NA2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211B100M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211B100M1R (A1, B, C, NA2, Z);
  input A1, B, C, NA2;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(B_bar, B);
    buf SMC_I3(OUT1, B_bar);
    not SMC_I4(A1_bar, A1);
    and SMC_I5(OUT2, A1_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && C===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && C===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && C===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && B===1'b1 && NA2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && B===1'b1 && NA2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && B===1'b1 && NA2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211B100M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211B100M2R (A1, B, C, NA2, Z);
  input A1, B, C, NA2;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(B_bar, B);
    buf SMC_I3(OUT1, B_bar);
    not SMC_I4(A1_bar, A1);
    and SMC_I5(OUT2, A1_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && C===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && C===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && C===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && B===1'b1 && NA2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && B===1'b1 && NA2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && B===1'b1 && NA2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211B100M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211B100M4R (A1, B, C, NA2, Z);
  input A1, B, C, NA2;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(B_bar, B);
    buf SMC_I3(OUT1, B_bar);
    not SMC_I4(A1_bar, A1);
    and SMC_I5(OUT2, A1_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && C===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && C===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && C===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && B===1'b1 && NA2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && B===1'b1 && NA2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && B===1'b1 && NA2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211B100M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211B100M8RA (A1, B, C, NA2, Z);
  input A1, B, C, NA2;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(B_bar, B);
    buf SMC_I3(OUT1, B_bar);
    not SMC_I4(A1_bar, A1);
    and SMC_I5(OUT2, A1_bar, NA2);
    or SMC_I6(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && C===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && C===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && C===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && B===1'b1 && NA2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && B===1'b1 && NA2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && B===1'b1 && NA2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211B100M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211M0R (A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(A1_bar, A1);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A1_bar, A2_bar);
    not SMC_I5(B_bar, B);
    buf SMC_I6(OUT2, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211M1R (A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(A1_bar, A1);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A1_bar, A2_bar);
    not SMC_I5(B_bar, B);
    buf SMC_I6(OUT2, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211M2R (A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(A1_bar, A1);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A1_bar, A2_bar);
    not SMC_I5(B_bar, B);
    buf SMC_I6(OUT2, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211M4R (A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(A1_bar, A1);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A1_bar, A2_bar);
    not SMC_I5(B_bar, B);
    buf SMC_I6(OUT2, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211M6RA (A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(A1_bar, A1);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A1_bar, A2_bar);
    not SMC_I5(B_bar, B);
    buf SMC_I6(OUT2, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI211M8RA (A1, A2, B, C, Z);
  input A1, A2, B, C;
  output Z;

    not SMC_I0(C_bar, C);
    buf SMC_I1(OUT0, C_bar);
    not SMC_I2(A1_bar, A1);
    not SMC_I3(A2_bar, A2);
    and SMC_I4(OUT1, A1_bar, A2_bar);
    not SMC_I5(B_bar, B);
    buf SMC_I6(OUT2, B_bar);
    or SMC_I7(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI211M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M0R (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M12RA (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M16RA (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M1R (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M2R (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M4R (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M6RA (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B01M8RA (A1, A2, NB, Z);
  input A1, A2, NB;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    buf SMC_I3(OUT1, NB);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc NB --> Z
    if (A1===1'b0 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (NB => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (NB => Z) = (0.0, 0.0);
    ifnone
        (NB => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B01M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M0R (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M12RA (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M16RA (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M1R (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M2R (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M4R (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M6RA (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B10M8RA (A1, B, NA2, Z);
  input A1, B, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    not SMC_I2(A1_bar, A1);
    and SMC_I3(OUT1, A1_bar, NA2);
    or SMC_I4(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B10M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M0R (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M12RA (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M1R (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M2R (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M4R (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M6RA (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21B20M8RA (B, NA1, NA2, Z);
  input B, NA1, NA2;
  output Z;

    not SMC_I0(B_bar, B);
    buf SMC_I1(OUT0, B_bar);
    and SMC_I2(OUT1, NA1, NA2);
    or SMC_I3(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B --> Z
    if (NA1===1'b0 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b0 && NA2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (NA1===1'b1 && NA2===1'b0)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21B20M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M0R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M12RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M16RA (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M1R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M2R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M3R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M3R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M4R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M6R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI21M8R (A1, A2, B, Z);
  input A1, A2, B;
  output Z;

    not SMC_I0(A1_bar, A1);
    not SMC_I1(A2_bar, A2);
    and SMC_I2(OUT0, A1_bar, A2_bar);
    not SMC_I3(B_bar, B);
    buf SMC_I4(OUT1, B_bar);
    or SMC_I5(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI21M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI221M0R ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    or (tmp1, A1, A2);
    or (tmp2, B1, B2);
  nand (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI221M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI221M1R ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    or (tmp1, A1, A2);
    or (tmp2, B1, B2);
  nand (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI221M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI221M2R ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    or (tmp1, A1, A2);
    or (tmp2, B1, B2);
  nand (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI221M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI221M4R ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    or (tmp1, A1, A2);
    or (tmp2, B1, B2);
  nand (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI221M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI221M6RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    or (tmp1, A1, A2);
    or (tmp2, B1, B2);
  nand (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI221M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI221M8RA ( Z, A1, A2, B1, B2, C );
   input A1, A2, B1, B2, C;
   output Z;

    or (tmp1, A1, A2);
    or (tmp2, B1, B2);
  nand (Z, tmp1, tmp2, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI221M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI222M0RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

     or (tmp1, A1, A2);
     or (tmp2, B1, B2);
     or (tmp3, C1, C2);
   nand (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI222M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI222M1RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

     or (tmp1, A1, A2);
     or (tmp2, B1, B2);
     or (tmp3, C1, C2);
   nand (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI222M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI222M2RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

     or (tmp1, A1, A2);
     or (tmp2, B1, B2);
     or (tmp3, C1, C2);
   nand (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI222M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI222M4R ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

     or (tmp1, A1, A2);
     or (tmp2, B1, B2);
     or (tmp3, C1, C2);
   nand (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI222M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI222M6RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

     or (tmp1, A1, A2);
     or (tmp2, B1, B2);
     or (tmp3, C1, C2);
   nand (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI222M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI222M8RA ( Z, A1, A2, B1, B2, C1, C2 );
   input A1, A2, B1, B2, C1, C2;
   output Z;

     or (tmp1, A1, A2);
     or (tmp2, B1, B2);
     or (tmp3, C1, C2);
   nand (Z, tmp1, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b1 && C2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b0 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0 && C1===1'b1 && C2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b0 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && C1===1'b1 && C2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc C1 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C2===1'b0)
        (C1 => Z) = (0.0, 0.0);
    ifnone
        (C1 => Z) = (0.0, 0.0);

    // arc C2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b0 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b1 && B2===1'b1 && C1===1'b0)
        (C2 => Z) = (0.0, 0.0);
    ifnone
        (C2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI222M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22B10M0R ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;

    not (tmp1, NA2);
     or (tmp2, A1, tmp1);
     or (tmp3, B1, B2);
   nand (Z, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && B2===1'b1 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && B2===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && B1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B10M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22B10M1R ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;

    not (tmp1, NA2);
     or (tmp2, A1, tmp1);
     or (tmp3, B1, B2);
   nand (Z, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && B2===1'b1 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && B2===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && B1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B10M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22B10M2R ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;

    not (tmp1, NA2);
     or (tmp2, A1, tmp1);
     or (tmp3, B1, B2);
   nand (Z, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && B2===1'b1 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && B2===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && B1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B10M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22B10M4R ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;

    not (tmp1, NA2);
     or (tmp2, A1, tmp1);
     or (tmp3, B1, B2);
   nand (Z, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && B2===1'b1 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && B2===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && B1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B10M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22B10M8RA ( Z, A1, B1, B2, NA2 );
   input A1, B1, B2, NA2;
   output Z;

    not (tmp1, NA2);
     or (tmp2, A1, tmp1);
     or (tmp3, B1, B2);
   nand (Z, tmp2, tmp3);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (B1===1'b0 && B2===1'b1 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && B2===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B2===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && B1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && B1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (NA2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B10M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22B20M0R ( Z, B1, B2, NA1, NA2 );
   input B1, B2, NA1, NA2;
   output Z;

     nand (tmp1, NA1, NA2);
       or (tmp2, B1,  B2);
     nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    if (B2===1'b0 && NA1===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b0 && NA1===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b0 && NA1===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (B1===1'b0 && NA1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    if (B1===1'b0 && B2===1'b1 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    ifnone
        (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (B1===1'b0 && B2===1'b1 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B20M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22B20M1R ( Z, B1, B2, NA1, NA2 );
   input B1, B2, NA1, NA2;
   output Z;

     nand (tmp1, NA1, NA2);
       or (tmp2, B1,  B2);
     nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    if (B2===1'b0 && NA1===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b0 && NA1===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b0 && NA1===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (B1===1'b0 && NA1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    if (B1===1'b0 && B2===1'b1 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    ifnone
        (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (B1===1'b0 && B2===1'b1 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B20M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22B20M2R ( Z, B1, B2, NA1, NA2 );
   input B1, B2, NA1, NA2;
   output Z;

     nand (tmp1, NA1, NA2);
       or (tmp2, B1,  B2);
     nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    if (B2===1'b0 && NA1===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b0 && NA1===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b0 && NA1===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (B1===1'b0 && NA1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    if (B1===1'b0 && B2===1'b1 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    ifnone
        (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (B1===1'b0 && B2===1'b1 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B20M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22B20M4R ( Z, B1, B2, NA1, NA2 );
   input B1, B2, NA1, NA2;
   output Z;

     nand (tmp1, NA1, NA2);
       or (tmp2, B1,  B2);
     nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    if (B2===1'b0 && NA1===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b0 && NA1===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b0 && NA1===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (B1===1'b0 && NA1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    if (B1===1'b0 && B2===1'b1 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    ifnone
        (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (B1===1'b0 && B2===1'b1 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B20M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22B20M8RA ( Z, B1, B2, NA1, NA2 );
   input B1, B2, NA1, NA2;
   output Z;

     nand (tmp1, NA1, NA2);
       or (tmp2, B1,  B2);
     nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc B1 --> Z
    if (B2===1'b0 && NA1===1'b0 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b0 && NA1===1'b0 && NA2===1'b1)
        (B1 => Z) = (0.0, 0.0);
    if (B2===1'b0 && NA1===1'b1 && NA2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (B1===1'b0 && NA1===1'b0 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA1===1'b0 && NA2===1'b1)
        (B2 => Z) = (0.0, 0.0);
    if (B1===1'b0 && NA1===1'b1 && NA2===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc NA1 --> Z
    if (B1===1'b0 && B2===1'b1 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA2===1'b1)
        (NA1 => Z) = (0.0, 0.0);
    ifnone
        (NA1 => Z) = (0.0, 0.0);

    // arc NA2 --> Z
    if (B1===1'b0 && B2===1'b1 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b0 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    if (B1===1'b1 && B2===1'b1 && NA1===1'b1)
        (NA2 => Z) = (0.0, 0.0);
    ifnone
        (NA2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22B20M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22M0R ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

      or (tmp1, A1, A2);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22M12RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

      or (tmp1, A1, A2);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22M16RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

      or (tmp1, A1, A2);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22M1R ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

      or (tmp1, A1, A2);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22M2R ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

      or (tmp1, A1, A2);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22M4R ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

      or (tmp1, A1, A2);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22M6RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

      or (tmp1, A1, A2);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI22M8RA ( Z, A1, A2, B1, B2 );
   input A1, A2, B1, B2;
   output Z;

      or (tmp1, A1, A2);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI22M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI31M0R ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;

    or (tmp1, A1, A2, A3);
  nand (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI31M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI31M1R ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;

    or (tmp1, A1, A2, A3);
  nand (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI31M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI31M2R ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;

    or (tmp1, A1, A2, A3);
  nand (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI31M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI31M4R ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;

    or (tmp1, A1, A2, A3);
  nand (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI31M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI31M8RA ( Z, A1, A2, A3, B );
   input A1, A2, A3, B;
   output Z;

    or (tmp1, A1, A2, A3);
  nand (Z, tmp1, B);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    (A3 => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI31M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI32M0R ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;

      or (tmp1, A1, A2, A3);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI32M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI32M1R ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;

      or (tmp1, A1, A2, A3);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI32M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI32M2R ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;

      or (tmp1, A1, A2, A3);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI32M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI32M4R ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;

      or (tmp1, A1, A2, A3);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI32M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI32M8RA ( Z, A1, A2, A3, B1, B2 );
   input A1, A2, A3, B1, B2;
   output Z;

      or (tmp1, A1, A2, A3);
      or (tmp2, B1, B2);
    nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI32M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI33M0R ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;

    or (tmp1, A1, A2, A3);
    or (tmp2, B1, B2, B3);
  nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI33M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI33M1R ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;

    or (tmp1, A1, A2, A3);
    or (tmp2, B1, B2, B3);
  nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI33M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI33M2R ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;

    or (tmp1, A1, A2, A3);
    or (tmp2, B1, B2, B3);
  nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI33M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI33M4R ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;

    or (tmp1, A1, A2, A3);
    or (tmp2, B1, B2, B3);
  nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI33M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OAI33M8RA ( Z, A1, A2, A3, B1, B2, B3 );
   input A1, A2, A3, B1, B2, B3;
   output Z;

    or (tmp1, A1, A2, A3);
    or (tmp2, B1, B2, B3);
  nand (Z, tmp1, tmp2);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A1 --> Z
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A1 => Z) = (0.0, 0.0);
    if (A2===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A1 => Z) = (0.0, 0.0);
    ifnone
        (A1 => Z) = (0.0, 0.0);

    // arc A2 --> Z
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A3===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A2 => Z) = (0.0, 0.0);
    ifnone
        (A2 => Z) = (0.0, 0.0);

    // arc A3 --> Z
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b0 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b0 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b0)
        (A3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b0 && B1===1'b1 && B2===1'b1 && B3===1'b1)
        (A3 => Z) = (0.0, 0.0);
    ifnone
        (A3 => Z) = (0.0, 0.0);

    // arc B1 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B2===1'b0 && B3===1'b0)
        (B1 => Z) = (0.0, 0.0);
    ifnone
        (B1 => Z) = (0.0, 0.0);

    // arc B2 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B3===1'b0)
        (B2 => Z) = (0.0, 0.0);
    ifnone
        (B2 => Z) = (0.0, 0.0);

    // arc B3 --> Z
    if (A1===1'b0 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b0 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b0 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b0 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    if (A1===1'b1 && A2===1'b1 && A3===1'b1 && B1===1'b0 && B2===1'b0)
        (B3 => Z) = (0.0, 0.0);
    ifnone
        (B3 => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OAI33M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M0R (A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR2M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M12RA (A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR2M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M16RA (A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR2M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M1R (A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR2M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M22RA (A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR2M22RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M2R (A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR2M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M4R (A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR2M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M6R (A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR2M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR2M8R (A, B, Z);
  input A, B;
  output Z;

    buf SMC_I0(OUT0, A);
    buf SMC_I1(OUT1, B);
    or SMC_I2(Z, OUT0, OUT1);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR2M8R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M0R (A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR3M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M12RA (A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR3M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M16RA (A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR3M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M1R (A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR3M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M2R (A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR3M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M4R (A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR3M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M6R (A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR3M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR3M8RA (A, B, C, Z);
  input A, B, C;
  output Z;

    buf SMC_I0(OUT0, B);
    buf SMC_I1(OUT1, A);
    buf SMC_I2(OUT2, C);
    or SMC_I3(Z, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR3M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M0R (A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR4M0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M12RA (A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR4M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M16RA (A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR4M16RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M1R (A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR4M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M2R (A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR4M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M4RA (A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR4M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M6R (A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR4M6R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR4M8RA (A, B, C, D, Z);
  input A, B, C, D;
  output Z;

    buf SMC_I0(OUT0, D);
    buf SMC_I1(OUT1, B);
    buf SMC_I2(OUT2, C);
    buf SMC_I3(OUT3, A);
    or SMC_I4(Z, OUT0, OUT1, OUT2, OUT3);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR4M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR6M12RA (A, B, C, D, E, F, Z);
  input A, B, C, D, E, F;
  output Z;

    buf SMC_I0(OUT0, F);
    buf SMC_I1(OUT1, C);
    buf SMC_I2(OUT2, A);
    buf SMC_I3(OUT3, B);
    buf SMC_I4(OUT4, D);
    buf SMC_I5(OUT5, E);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0, 0.0);

    // arc F --> Z
    (F => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR6M12RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR6M1RA (A, B, C, D, E, F, Z);
  input A, B, C, D, E, F;
  output Z;

    buf SMC_I0(OUT0, F);
    buf SMC_I1(OUT1, C);
    buf SMC_I2(OUT2, A);
    buf SMC_I3(OUT3, B);
    buf SMC_I4(OUT4, D);
    buf SMC_I5(OUT5, E);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0, 0.0);

    // arc F --> Z
    (F => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR6M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR6M2RA (A, B, C, D, E, F, Z);
  input A, B, C, D, E, F;
  output Z;

    buf SMC_I0(OUT0, F);
    buf SMC_I1(OUT1, C);
    buf SMC_I2(OUT2, A);
    buf SMC_I3(OUT3, B);
    buf SMC_I4(OUT4, D);
    buf SMC_I5(OUT5, E);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0, 0.0);

    // arc F --> Z
    (F => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR6M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR6M4RA (A, B, C, D, E, F, Z);
  input A, B, C, D, E, F;
  output Z;

    buf SMC_I0(OUT0, F);
    buf SMC_I1(OUT1, C);
    buf SMC_I2(OUT2, A);
    buf SMC_I3(OUT3, B);
    buf SMC_I4(OUT4, D);
    buf SMC_I5(OUT5, E);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0, 0.0);

    // arc F --> Z
    (F => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR6M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR6M6RA (A, B, C, D, E, F, Z);
  input A, B, C, D, E, F;
  output Z;

    buf SMC_I0(OUT0, F);
    buf SMC_I1(OUT1, C);
    buf SMC_I2(OUT2, A);
    buf SMC_I3(OUT3, B);
    buf SMC_I4(OUT4, D);
    buf SMC_I5(OUT5, E);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0, 0.0);

    // arc F --> Z
    (F => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR6M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module OR6M8RA (A, B, C, D, E, F, Z);
  input A, B, C, D, E, F;
  output Z;

    buf SMC_I0(OUT0, F);
    buf SMC_I1(OUT1, C);
    buf SMC_I2(OUT2, A);
    buf SMC_I3(OUT3, B);
    buf SMC_I4(OUT4, D);
    buf SMC_I5(OUT5, E);
    or SMC_I6(Z, OUT0, OUT1, OUT2, OUT3, OUT4, OUT5);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    (A => Z) = (0.0, 0.0);

    // arc B --> Z
    (B => Z) = (0.0, 0.0);

    // arc C --> Z
    (C => Z) = (0.0, 0.0);

    // arc D --> Z
    (D => Z) = (0.0, 0.0);

    // arc E --> Z
    (E => Z) = (0.0, 0.0);

    // arc F --> Z
    (F => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // OR6M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module REG1M1R (RD, RG, RGB, WE, RQB);
  input RD, RG, RGB, WE;
  output RQB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(RD), .en(WE), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I1(.q(SMC_IQ), .d(RD), .en(WE), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(SMC_DINRQB, SMC_IQN);

    not SMC_I3(RGB_bar, RGB);
    nand SMC_I4(SMC_ZENRQB, RG, RGB_bar);


    bufif0 SMC_I5(RQB, SMC_DINRQB, SMC_ZENRQB);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I6(shcheckWERDhl, RG, RGB_bar);


  specify


    // arc RD --> RQB
    (RD => RQB) = (0.0, 0.0);

    // arc RG --> RQB
    if (RD===1'b0 && RGB===1'b0 && WE===1'b0)
    	(RG => RQB) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b0 && RGB===1'b0 && WE===1'b1)
    	(RG => RQB) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RGB===1'b0 && WE===1'b1)
    	(RG => RQB) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RGB===1'b0 && WE===1'b0)
    	(RG => RQB) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    ifnone
    	(RG => RQB) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);

    // arc RGB --> RQB
    if (RD===1'b1 && RG===1'b1 && WE===1'b1)
    	(RGB => RQB) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b0 && RG===1'b1 && WE===1'b1)
    	(RGB => RQB) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RG===1'b1 && WE===1'b0)
    	(RGB => RQB) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b0 && RG===1'b1 && WE===1'b0)
    	(RGB => RQB) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    ifnone
    	(RGB => RQB) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);

    // arc WE --> RQB
    (posedge WE => ( RQB +: RD )) = (0.0, 0.0);



    // setup
    $setup( negedge RD, negedge WE &&&
        (shcheckWERDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RD, negedge WE &&&
        (shcheckWERDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge WE &&&
        (shcheckWERDhl === 1'b1), negedge RD, 0.0, notifier );

    // hold
    $hold( negedge WE &&&
        (shcheckWERDhl === 1'b1), posedge RD, 0.0, notifier );

    // mpw
    $width( posedge WE, 0.0, 0, notifier );

    // mpw
    $width( negedge WE, 0.0, 0, notifier );

    $period( posedge WE, 0, notifier );
    $period( negedge WE, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // REG1M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module REG2M1R (RD, RG1, RG2, WE, RQ1B, RQ2B);
  input RD, RG1, RG2, WE;
  output RQ1B, RQ2B;
  reg notifier;

  wire SMC_LD_IN;
    not SMC_I0(SMC_LD_IN, RD);

    not SMC_I1(SMC_IQN, SMC_IQ);

  `ifdef functional // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(SMC_LD_IN), .en(WE), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    ldlatch_p0 SMC_I2(.q(SMC_IQ), .d(SMC_LD_IN), .en(WE), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(SMC_DINRQ1B, SMC_IQ);

    not SMC_I4(SMC_ZENRQ1B, RG1);


    bufif0 SMC_I5(RQ1B, SMC_DINRQ1B, SMC_ZENRQ1B);

    buf SMC_I6(SMC_DINRQ2B, SMC_IQ);

    not SMC_I7(SMC_ZENRQ2B, RG2);


    bufif0 SMC_I8(RQ2B, SMC_DINRQ2B, SMC_ZENRQ2B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc RD --> RQ1B
    if (RG1===1'b1 && RG2===1'b0 && WE===1'b1)
        (RD => RQ1B) = (0.0, 0.0);
    if (RG1===1'b1 && RG2===1'b1 && WE===1'b1)
        (RD => RQ1B) = (0.0, 0.0);
    ifnone
    	(RD => RQ1B) = (0.0, 0.0);

    // arc RD --> RQ2B
    if (RG1===1'b0 && RG2===1'b1 && WE===1'b1)
        (RD => RQ2B) = (0.0, 0.0);
    if (RG1===1'b1 && RG2===1'b1 && WE===1'b1)
        (RD => RQ2B) = (0.0, 0.0);
    ifnone
    	(RD => RQ2B) = (0.0, 0.0);

    // arc RG1 --> RQ1B
    if (RD===1'b0 && RG2===1'b0 && WE===1'b0)
    	(RG1 => RQ1B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b0 && RG2===1'b1 && WE===1'b0)
    	(RG1 => RQ1B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RG2===1'b0 && WE===1'b0)
    	(RG1 => RQ1B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RG2===1'b1 && WE===1'b0)
    	(RG1 => RQ1B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b0 && RG2===1'b0 && WE===1'b1)
    	(RG1 => RQ1B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b0 && RG2===1'b1 && WE===1'b1)
    	(RG1 => RQ1B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RG2===1'b0 && WE===1'b1)
    	(RG1 => RQ1B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RG2===1'b1 && WE===1'b1)
    	(RG1 => RQ1B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    ifnone
    	(RG1 => RQ1B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);

    // arc RG2 --> RQ2B
    if (RD===1'b0 && RG1===1'b0 && WE===1'b0)
    	(RG2 => RQ2B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b0 && RG1===1'b1 && WE===1'b0)
    	(RG2 => RQ2B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RG1===1'b0 && WE===1'b0)
    	(RG2 => RQ2B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RG1===1'b1 && WE===1'b0)
    	(RG2 => RQ2B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b0 && RG1===1'b0 && WE===1'b1)
    	(RG2 => RQ2B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b0 && RG1===1'b1 && WE===1'b1)
    	(RG2 => RQ2B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RG1===1'b0 && WE===1'b1)
    	(RG2 => RQ2B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    if (RD===1'b1 && RG1===1'b1 && WE===1'b1)
    	(RG2 => RQ2B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);
    ifnone
    	(RG2 => RQ1B) = (0.0, 0.0, 0.0, 0.0, 0.0, 0.0);

    // arc WE --> RQ1B
    if (RD===1'b1 && RG1===1'b1 && RG2===1'b0)
    	(posedge WE => ( RQ1B -: RD )) = (0.0, 0.0);
    if (RD===1'b0 && RG1===1'b1 && RG2===1'b0)
    	(posedge WE => ( RQ1B -: RD )) = (0.0, 0.0);
    if (RD===1'b1 && RG1===1'b1 && RG2===1'b1)
    	(posedge WE => ( RQ1B -: RD )) = (0.0, 0.0);
    if (RD===1'b0 && RG1===1'b1 && RG2===1'b1)
    	(posedge WE => ( RQ1B -: RD )) = (0.0, 0.0);
    ifnone
    	(posedge WE => ( RQ1B -: RD )) = (0.0, 0.0);

    // arc WE --> RQ2B
    if (RD===1'b1 && RG1===1'b0 && RG2===1'b1)
    	(posedge WE => ( RQ2B -: RD )) = (0.0, 0.0);
    if (RD===1'b0 && RG1===1'b0 && RG2===1'b1)
    	(posedge WE => ( RQ2B -: RD )) = (0.0, 0.0);
    if (RD===1'b1 && RG1===1'b1 && RG2===1'b1)
    	(posedge WE => ( RQ2B -: RD )) = (0.0, 0.0);
    if (RD===1'b0 && RG1===1'b1 && RG2===1'b1)
    	(posedge WE => ( RQ2B -: RD )) = (0.0, 0.0);
    ifnone
    	(posedge WE => ( RQ2B -: RD )) = (0.0, 0.0);



    // setup
    $setup( posedge RD, negedge WE, 0.0, notifier );

    // setup
    $setup( negedge RD, negedge WE, 0.0, notifier );

    // hold
    $hold( negedge WE, posedge RD, 0.0, notifier );

    // hold
    $hold( negedge WE, negedge RD, 0.0, notifier );

    // mpw
    $width( posedge WE, 0.0, 0, notifier );

    // mpw
    $width( negedge WE, 0.0, 0, notifier );

    $period( posedge WE, 0, notifier );
    $period( negedge WE, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // REG2M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module REGKM1R (RD, RQB);
  input RD;
  output RQB;
  reg NOTIFIER;

    buf(weak0,weak1) SMC_IO(RD, io_wire);
    buf              SMC_I1(io_wire, RD);
    not              SMC_I0(RQB, RD);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc RD --> RQB
    (RD => RQB) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // REGKM1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module REGKM2R (RD, RQB);
  input RD;
  output RQB;
  reg NOTIFIER;

    buf(weak0,weak1) SMC_IO(RD, io_wire);
    buf              SMC_I1(io_wire, RD);
    not              SMC_I0(RQB, RD);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc RD --> RQB
    (RD => RQB) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // REGKM2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module REGKM4R (RD, RQB);
  input RD;
  output RQB;
  reg NOTIFIER;

    buf(weak0,weak1) SMC_IO(RD, io_wire);
    buf              SMC_I1(io_wire, RD);
    not              SMC_I0(RQB, RD);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc RD --> RQB
    (RD => RQB) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // REGKM4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFAQM1RA (A, B, SD, SE, CK, Q);
  input A, B, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, A, B, SE_bar);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKAlh, SE);

    not SMC_I7(shcheckCKBlh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: B )) = (0.0, 0.0);



    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge B, posedge CK &&&
        (shcheckCKBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge B, posedge CK &&&
        (shcheckCKBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge A, posedge CK &&&
        (shcheckCKAlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge A, posedge CK &&&
        (shcheckCKAlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKBlh === 1'b1), posedge B, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKBlh === 1'b1), negedge B, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKAlh === 1'b1), posedge A, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKAlh === 1'b1), negedge A, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFAQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFAQM2RA (A, B, SD, SE, CK, Q);
  input A, B, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, A, B, SE_bar);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKAlh, SE);

    not SMC_I7(shcheckCKBlh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: B )) = (0.0, 0.0);



    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge B, posedge CK &&&
        (shcheckCKBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge B, posedge CK &&&
        (shcheckCKBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge A, posedge CK &&&
        (shcheckCKAlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge A, posedge CK &&&
        (shcheckCKAlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKBlh === 1'b1), posedge B, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKBlh === 1'b1), negedge B, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKAlh === 1'b1), posedge A, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKAlh === 1'b1), negedge A, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFAQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFAQM4RA (A, B, SD, SE, CK, Q);
  input A, B, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, A, B, SE_bar);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKAlh, SE);

    not SMC_I7(shcheckCKBlh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: B )) = (0.0, 0.0);



    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge B, posedge CK &&&
        (shcheckCKBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge B, posedge CK &&&
        (shcheckCKBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge A, posedge CK &&&
        (shcheckCKAlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge A, posedge CK &&&
        (shcheckCKAlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKBlh === 1'b1), posedge B, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKBlh === 1'b1), negedge B, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKAlh === 1'b1), posedge A, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKAlh === 1'b1), negedge A, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFAQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFAQM6RA (A, B, SD, SE, CK, Q);
  input A, B, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, A, B, SE_bar);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKAlh, SE);

    not SMC_I7(shcheckCKBlh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: B )) = (0.0, 0.0);



    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge B, posedge CK &&&
        (shcheckCKBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge B, posedge CK &&&
        (shcheckCKBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge A, posedge CK &&&
        (shcheckCKAlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge A, posedge CK &&&
        (shcheckCKAlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKBlh === 1'b1), posedge B, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKBlh === 1'b1), negedge B, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKAlh === 1'b1), posedge A, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKAlh === 1'b1), negedge A, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFAQM6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFAQM8RA (A, B, SD, SE, CK, Q);
  input A, B, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, A, B, SE_bar);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKAlh, SE);

    not SMC_I7(shcheckCKBlh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: B )) = (0.0, 0.0);



    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge B, posedge CK &&&
        (shcheckCKBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge B, posedge CK &&&
        (shcheckCKBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge A, posedge CK &&&
        (shcheckCKAlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge A, posedge CK &&&
        (shcheckCKAlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKBlh === 1'b1), posedge B, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKBlh === 1'b1), negedge B, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKAlh === 1'b1), posedge A, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKAlh === 1'b1), negedge A, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFAQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCM1RA (D, SD, SE, CKB, Q, QB);
  input D, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKBDhl, SE);

    buf SMC_I7(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CKB-lh (!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // setup D-lh CKB-lh (!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // setup SE-hl CKB-lh ()
    $setup(negedge SE, negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-lh ()
    $setup(posedge SE, negedge CKB, 0.0, notifier);

    // setup SD-hl CKB-lh (SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // setup SD-lh CKB-lh (SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // hold D-hl CKB-lh (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // hold D-lh CKB-lh (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // hold SE-hl CKB-lh ()
    $hold(negedge CKB, negedge SE, 0.0, notifier);

    // hold SE-lh CKB-lh ()
    $hold(negedge CKB, posedge SE, 0.0, notifier);

    // hold SD-hl CKB-lh (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // hold SD-lh CKB-lh (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(posedge CKB, 0.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(negedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCM2RA (D, SD, SE, CKB, Q, QB);
  input D, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKBDhl, SE);

    buf SMC_I7(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CKB-lh (!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // setup D-lh CKB-lh (!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // setup SE-hl CKB-lh ()
    $setup(negedge SE, negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-lh ()
    $setup(posedge SE, negedge CKB, 0.0, notifier);

    // setup SD-hl CKB-lh (SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // setup SD-lh CKB-lh (SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // hold D-hl CKB-lh (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // hold D-lh CKB-lh (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // hold SE-hl CKB-lh ()
    $hold(negedge CKB, negedge SE, 0.0, notifier);

    // hold SE-lh CKB-lh ()
    $hold(negedge CKB, posedge SE, 0.0, notifier);

    // hold SD-hl CKB-lh (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // hold SD-lh CKB-lh (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(posedge CKB, 0.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(negedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCM4RA (D, SD, SE, CKB, Q, QB);
  input D, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKBDhl, SE);

    buf SMC_I7(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CKB-lh (!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // setup D-lh CKB-lh (!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // setup SE-hl CKB-lh ()
    $setup(negedge SE, negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-lh ()
    $setup(posedge SE, negedge CKB, 0.0, notifier);

    // setup SD-hl CKB-lh (SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // setup SD-lh CKB-lh (SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // hold D-hl CKB-lh (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // hold D-lh CKB-lh (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // hold SE-hl CKB-lh ()
    $hold(negedge CKB, negedge SE, 0.0, notifier);

    // hold SE-lh CKB-lh ()
    $hold(negedge CKB, posedge SE, 0.0, notifier);

    // hold SD-hl CKB-lh (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // hold SD-lh CKB-lh (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(posedge CKB, 0.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(negedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCM8RA (D, SD, SE, CKB, Q, QB);
  input D, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKBDhl, SE);

    buf SMC_I7(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge CKB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CKB-lh (!SE)
    $setup(negedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // setup D-lh CKB-lh (!SE)
    $setup(posedge D &&& (shcheckCKBDhl === 1'b1),
        negedge CKB &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // setup SE-hl CKB-lh ()
    $setup(negedge SE, negedge CKB, 0.0, notifier);

    // setup SE-lh CKB-lh ()
    $setup(posedge SE, negedge CKB, 0.0, notifier);

    // setup SD-hl CKB-lh (SE)
    $setup(negedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // setup SD-lh CKB-lh (SE)
    $setup(posedge SD &&& (shcheckCKBSDhl === 1'b1),
        negedge CKB &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // hold D-hl CKB-lh (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        negedge D &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // hold D-lh CKB-lh (!SE)
    $hold(negedge CKB &&& (shcheckCKBDhl === 1'b1),
        posedge D &&& (shcheckCKBDhl === 1'b1), 0.0, notifier);

    // hold SE-hl CKB-lh ()
    $hold(negedge CKB, negedge SE, 0.0, notifier);

    // hold SE-lh CKB-lh ()
    $hold(negedge CKB, posedge SE, 0.0, notifier);

    // hold SD-hl CKB-lh (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        negedge SD &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // hold SD-lh CKB-lh (SE)
    $hold(negedge CKB &&& (shcheckCKBSDhl === 1'b1),
        posedge SD &&& (shcheckCKBSDhl === 1'b1), 0.0, notifier);

    // mpw CKB-hl NS-hl ()
    $width(posedge CKB, 0.0, 0, notifier);

    // mpw CKB-lh NS-lh ()
    $width(negedge CKB, 0.0, 0, notifier);

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQM1RA (D, SD, SE, CKB, Q);
  input D, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKBDhl, SE);

    buf SMC_I5(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB, 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB, 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB, negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB, posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQM2RA (D, SD, SE, CKB, Q);
  input D, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKBDhl, SE);

    buf SMC_I5(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB, 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB, 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB, negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB, posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQM4RA (D, SD, SE, CKB, Q);
  input D, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKBDhl, SE);

    buf SMC_I5(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB, 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB, 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB, negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB, posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQM8RA (D, SD, SE, CKB, Q);
  input D, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKBDhl, SE);

    buf SMC_I5(shcheckCKBSDhl, SE);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB, 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB, 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB, negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB, posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQRM1RA (D, RB, SD, SE, CKB, Q);
  input D, RB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, RB, SE_bar);

    and SMC_I6(shcheckCKBSDhl, RB, SE);

    buf SMC_I7(shcheckCKBSEhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQRM2RA (D, RB, SD, SE, CKB, Q);
  input D, RB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, RB, SE_bar);

    and SMC_I6(shcheckCKBSDhl, RB, SE);

    buf SMC_I7(shcheckCKBSEhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQRM4RA (D, RB, SD, SE, CKB, Q);
  input D, RB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, RB, SE_bar);

    and SMC_I6(shcheckCKBSDhl, RB, SE);

    buf SMC_I7(shcheckCKBSEhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQRM8RA (D, RB, SD, SE, CKB, Q);
  input D, RB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, RB, SE_bar);

    and SMC_I6(shcheckCKBSDhl, RB, SE);

    buf SMC_I7(shcheckCKBSEhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQRSM1RA (D, RB, SB, SD, SE, CKB, Q);
  input D, RB, SB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKBRBhl, SB);

    buf SMC_I7(shcheckCKBSBhl, RB);

    and SMC_I8(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I9(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQRSM2RA (D, RB, SB, SD, SE, CKB, Q);
  input D, RB, SB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKBRBhl, SB);

    buf SMC_I7(shcheckCKBSBhl, RB);

    and SMC_I8(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I9(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQRSM4RA (D, RB, SB, SD, SE, CKB, Q);
  input D, RB, SB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKBRBhl, SB);

    buf SMC_I7(shcheckCKBSBhl, RB);

    and SMC_I8(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I9(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQRSM8RA (D, RB, SB, SD, SE, CKB, Q);
  input D, RB, SB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I6(shcheckCKBRBhl, SB);

    buf SMC_I7(shcheckCKBSBhl, RB);

    and SMC_I8(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I9(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQSM1RA (D, SB, SD, SE, CKB, Q);
  input D, SB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, SB, SE_bar);

    and SMC_I6(shcheckCKBSDhl, SB, SE);

    buf SMC_I7(shcheckCKBSEhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQSM2RA (D, SB, SD, SE, CKB, Q);
  input D, SB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, SB, SE_bar);

    and SMC_I6(shcheckCKBSDhl, SB, SE);

    buf SMC_I7(shcheckCKBSEhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQSM4RA (D, SB, SD, SE, CKB, Q);
  input D, SB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, SB, SE_bar);

    and SMC_I6(shcheckCKBSDhl, SB, SE);

    buf SMC_I7(shcheckCKBSEhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCQSM8RA (D, SB, SD, SE, CKB, Q);
  input D, SB, SD, SE, CKB;
  output Q;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKBDhl, SB, SE_bar);

    and SMC_I6(shcheckCKBSDhl, SB, SE);

    buf SMC_I7(shcheckCKBSEhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCQSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCRM1RA (D, RB, SD, SE, CKB, Q, QB);
  input D, RB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, RB, SE_bar);

    and SMC_I8(shcheckCKBSDhl, RB, SE);

    buf SMC_I9(shcheckCKBSEhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCRM2RA (D, RB, SD, SE, CKB, Q, QB);
  input D, RB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, RB, SE_bar);

    and SMC_I8(shcheckCKBSDhl, RB, SE);

    buf SMC_I9(shcheckCKBSEhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCRM4RA (D, RB, SD, SE, CKB, Q, QB);
  input D, RB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, RB, SE_bar);

    and SMC_I8(shcheckCKBSDhl, RB, SE);

    buf SMC_I9(shcheckCKBSEhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCRM8RA (D, RB, SD, SE, CKB, Q, QB);
  input D, RB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, RB, SE_bar);

    and SMC_I8(shcheckCKBSDhl, RB, SE);

    buf SMC_I9(shcheckCKBSEhl, RB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCRSM1RA (D, RB, SB, SD, SE, CKB, Q, QB);
  input D, RB, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I8(shcheckCKBRBhl, SB);

    buf SMC_I9(shcheckCKBSBhl, RB);

    and SMC_I10(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I11(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCRSM2RA (D, RB, SB, SD, SE, CKB, Q, QB);
  input D, RB, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I8(shcheckCKBRBhl, SB);

    buf SMC_I9(shcheckCKBSBhl, RB);

    and SMC_I10(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I11(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCRSM4RA (D, RB, SB, SD, SE, CKB, Q, QB);
  input D, RB, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I8(shcheckCKBRBhl, SB);

    buf SMC_I9(shcheckCKBSBhl, RB);

    and SMC_I10(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I11(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCRSM8RA (D, RB, SB, SD, SE, CKB, Q, QB);
  input D, RB, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);


    inv_clr0 SMC_I1(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB) );

  `else // functional //

    dff_p0 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(RB), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, RB, SB, SE_bar);

    buf SMC_I8(shcheckCKBRBhl, SB);

    buf SMC_I9(shcheckCKBSBhl, RB);

    and SMC_I10(shcheckCKBSDhl, RB, SB, SE);

    and SMC_I11(shcheckCKBSEhl, RB, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBRBhl === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( negedge CKB &&&
        (shcheckCKBSBhl === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCSM1RA (D, SB, SD, SE, CKB, Q, QB);
  input D, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB) );

  `else // functional //

    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, SB, SE_bar);

    and SMC_I8(shcheckCKBSDhl, SB, SE);

    buf SMC_I9(shcheckCKBSEhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCSM2RA (D, SB, SD, SE, CKB, Q, QB);
  input D, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB) );

  `else // functional //

    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, SB, SE_bar);

    and SMC_I8(shcheckCKBSDhl, SB, SE);

    buf SMC_I9(shcheckCKBSEhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCSM4RA (D, SB, SD, SE, CKB, Q, QB);
  input D, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB) );

  `else // functional //

    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, SB, SE_bar);

    and SMC_I8(shcheckCKBSDhl, SB, SE);

    buf SMC_I9(shcheckCKBSEhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFCSM8RA (D, SB, SD, SE, CKB, Q, QB);
  input D, SB, SD, SE, CKB;
  output Q, QB;
  reg notifier;

    wire SMC_CK_IN;
    not SMC_I0(SMC_CK_IN, CKB);

    not SMC_I1(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I2(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB) );

  `else // functional //

    dff_p1 SMC_I3(.q(SMC_IQ), .d(SMC_NS_IN), .clk(SMC_CK_IN),
          .clear(1'b1), .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I4(Q, SMC_IQ);

    buf SMC_I5(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(SE_bar, SE);
    and SMC_I7(shcheckCKBDhl, SB, SE_bar);

    and SMC_I8(shcheckCKBSDhl, SB, SE);

    buf SMC_I9(shcheckCKBSEhl, SB);


  specify


    // arc CKB --> Q
    (negedge CKB => ( Q +: D )) = (0.0, 0.0);

    // arc CKB --> QB
    (negedge CKB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, negedge CKB &&&
        (shcheckCKBDhl === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSEhl === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBDhl === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( negedge CKB &&&
        (shcheckCKBSDhl === 1'b1), posedge SD, 0.0, notifier );

    // recovery
    $recovery( posedge SB, negedge CKB, 0.0, notifier );

    // removal
    $hold( negedge CKB, posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CKB, 0.0, 0, notifier );

    // mpw
    $width( posedge CKB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    $period( posedge CKB, 0, notifier );
    $period( negedge CKB, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFCSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEM1RA (D, E, SD, SE, CK, Q, QB);
  input D, E, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFE_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, SE_bar);

    not SMC_I7(shcheckCKElh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEM2RA (D, E, SD, SE, CK, Q, QB);
  input D, E, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFE_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, SE_bar);

    not SMC_I7(shcheckCKElh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEM4RA (D, E, SD, SE, CK, Q, QB);
  input D, E, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFE_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, SE_bar);

    not SMC_I7(shcheckCKElh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEM8RA (D, E, SD, SE, CK, Q, QB);
  input D, E, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFE_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, SE_bar);

    not SMC_I7(shcheckCKElh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQBM1RA (D, E, SD, SE, CK, QB);
  input D, E, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEQB_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, E, SE_bar);

    not SMC_I6(shcheckCKElh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQBM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQBM2RA (D, E, SD, SE, CK, QB);
  input D, E, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEQB_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, E, SE_bar);

    not SMC_I6(shcheckCKElh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQBM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQBM4RA (D, E, SD, SE, CK, QB);
  input D, E, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEQB_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, E, SE_bar);

    not SMC_I6(shcheckCKElh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQBM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQBM8RA (D, E, SD, SE, CK, QB);
  input D, E, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEQB_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, E, SE_bar);

    not SMC_I6(shcheckCKElh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    if (D===1'b1 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQBM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQM0RA (D, E, SD, SE, CK, Q);
  input D, E, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQ_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, SE_bar);

    not SMC_I5(shcheckCKElh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQM0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQM1RA (D, E, SD, SE, CK, Q);
  input D, E, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQ_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, SE_bar);

    not SMC_I5(shcheckCKElh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQM2RA (D, E, SD, SE, CK, Q);
  input D, E, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQ_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, SE_bar);

    not SMC_I5(shcheckCKElh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQM4RA (D, E, SD, SE, CK, Q);
  input D, E, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQ_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, SE_bar);

    not SMC_I5(shcheckCKElh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQM8RA (D, E, SD, SE, CK, Q);
  input D, E, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQ_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, SE_bar);

    not SMC_I5(shcheckCKElh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQRM1RA (D, E, RB, SD, SE, CK, Q);
  input D, E, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I5(shcheckCKElh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQRM2RA (D, E, RB, SD, SE, CK, Q);
  input D, E, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I5(shcheckCKElh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQRM4RA (D, E, RB, SD, SE, CK, Q);
  input D, E, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I5(shcheckCKElh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQRM8RA (D, E, RB, SD, SE, CK, Q);
  input D, E, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I5(shcheckCKElh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQZRM1RA (D, E, RB, SD, SE, CK, Q);
  input D, E, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQZR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I5(shcheckCKElh, RB, SE_bar);

    not SMC_I6(shcheckCKRBlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQZRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQZRM2RA (D, E, RB, SD, SE, CK, Q);
  input D, E, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQZR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I5(shcheckCKElh, RB, SE_bar);

    not SMC_I6(shcheckCKRBlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQZRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQZRM4RA (D, E, RB, SD, SE, CK, Q);
  input D, E, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQZR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I5(shcheckCKElh, RB, SE_bar);

    not SMC_I6(shcheckCKRBlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQZRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEQZRM8RA (D, E, RB, SD, SE, CK, Q);
  input D, E, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    SDFEQZR_UDP__OUT__ SMC_I0(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I5(shcheckCKElh, RB, SE_bar);

    not SMC_I6(shcheckCKRBlh, SE);

    buf SMC_I7(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEQZRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFERM1RA (D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFER_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I7(shcheckCKElh, RB, SE_bar);

    and SMC_I8(shcheckCKSDlh, RB, SE);

    buf SMC_I9(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: E )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFERM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFERM2RA (D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFER_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I7(shcheckCKElh, RB, SE_bar);

    and SMC_I8(shcheckCKSDlh, RB, SE);

    buf SMC_I9(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: E )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFERM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFERM4RA (D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFER_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I7(shcheckCKElh, RB, SE_bar);

    and SMC_I8(shcheckCKSDlh, RB, SE);

    buf SMC_I9(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: E )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFERM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFERM8RA (D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFER_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I7(shcheckCKElh, RB, SE_bar);

    and SMC_I8(shcheckCKSDlh, RB, SE);

    buf SMC_I9(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: E )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: E )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: E )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: E )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge E, posedge CK &&&
        (shcheckCKElh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), posedge E, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKElh === 1'b1), negedge E, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK, 0.0, notifier );

    // removal
    $hold( posedge CK, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFERM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEZRM1RA (D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEZR_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I7(shcheckCKElh, RB, SE_bar);

    not SMC_I8(shcheckCKRBlh, SE);

    buf SMC_I9(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (RB&!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (RB&!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEZRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEZRM2RA (D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEZR_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I7(shcheckCKElh, RB, SE_bar);

    not SMC_I8(shcheckCKRBlh, SE);

    buf SMC_I9(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (RB&!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (RB&!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEZRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEZRM4RA (D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEZR_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I7(shcheckCKElh, RB, SE_bar);

    not SMC_I8(shcheckCKRBlh, SE);

    buf SMC_I9(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (RB&!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (RB&!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEZRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFEZRM8RA (D, E, RB, SD, SE, CK, Q, QB);
  input D, E, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    SDFEZR_UDP__OUT__ SMC_I1(SMC_NS_IN, D, E, SMC_IQ, RB, SD, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, E, RB, SE_bar);

    and SMC_I7(shcheckCKElh, RB, SE_bar);

    not SMC_I8(shcheckCKRBlh, SE);

    buf SMC_I9(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && E===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup E-hl CK-lh (RB&!SE)
    $setup(negedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup E-lh CK-lh (RB&!SE)
    $setup(posedge E &&& (shcheckCKElh === 1'b1),
        posedge CK &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (E&RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-hl CK-lh (E&RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold E-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        negedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold E-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKElh === 1'b1),
        posedge E &&& (shcheckCKElh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (E&RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFEZRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFM1RA (D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(shcheckCKDlh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFM2RA (D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(shcheckCKDlh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFM4RA (D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(shcheckCKDlh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFM8RA (D, SD, SE, CK, Q, QB);
  input D, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(shcheckCKDlh, SE);

    buf SMC_I6(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFMM1RA (D1, D2, S, SD, SE, CK, Q, QB);
  input D1, D2, S, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(S_bar, S);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT0, D2, S_bar, SE_bar);
    and SMC_I4(OUT1, D1, S, SE_bar);
    and SMC_I5(OUT2, SD, SE);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I10(shcheckCKD1lh, S, SE_bar);

    and SMC_I11(shcheckCKD2lh, S_bar, SE_bar);

    buf SMC_I12(shcheckCKSDlh, SE);

    not SMC_I13(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFMM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFMM2RA (D1, D2, S, SD, SE, CK, Q, QB);
  input D1, D2, S, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(S_bar, S);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT0, D2, S_bar, SE_bar);
    and SMC_I4(OUT1, D1, S, SE_bar);
    and SMC_I5(OUT2, SD, SE);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I10(shcheckCKD1lh, S, SE_bar);

    and SMC_I11(shcheckCKD2lh, S_bar, SE_bar);

    buf SMC_I12(shcheckCKSDlh, SE);

    not SMC_I13(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFMM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFMM4RA (D1, D2, S, SD, SE, CK, Q, QB);
  input D1, D2, S, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(S_bar, S);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT0, D2, S_bar, SE_bar);
    and SMC_I4(OUT1, D1, S, SE_bar);
    and SMC_I5(OUT2, SD, SE);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I10(shcheckCKD1lh, S, SE_bar);

    and SMC_I11(shcheckCKD2lh, S_bar, SE_bar);

    buf SMC_I12(shcheckCKSDlh, SE);

    not SMC_I13(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFMM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFMM8RA (D1, D2, S, SD, SE, CK, Q, QB);
  input D1, D2, S, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(S_bar, S);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT0, D2, S_bar, SE_bar);
    and SMC_I4(OUT1, D1, S, SE_bar);
    and SMC_I5(OUT2, SD, SE);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I10(shcheckCKD1lh, S, SE_bar);

    and SMC_I11(shcheckCKD2lh, S_bar, SE_bar);

    buf SMC_I12(shcheckCKSDlh, SE);

    not SMC_I13(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFMM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFMQM1RA (D1, D2, S, SD, SE, CK, Q);
  input D1, D2, S, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(S_bar, S);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT0, D2, S_bar, SE_bar);
    and SMC_I3(OUT1, D1, S, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I8(shcheckCKD1lh, S, SE_bar);

    and SMC_I9(shcheckCKD2lh, S_bar, SE_bar);

    buf SMC_I10(shcheckCKSDlh, SE);

    not SMC_I11(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFMQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFMQM2RA (D1, D2, S, SD, SE, CK, Q);
  input D1, D2, S, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(S_bar, S);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT0, D2, S_bar, SE_bar);
    and SMC_I3(OUT1, D1, S, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I8(shcheckCKD1lh, S, SE_bar);

    and SMC_I9(shcheckCKD2lh, S_bar, SE_bar);

    buf SMC_I10(shcheckCKSDlh, SE);

    not SMC_I11(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFMQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFMQM4RA (D1, D2, S, SD, SE, CK, Q);
  input D1, D2, S, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(S_bar, S);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT0, D2, S_bar, SE_bar);
    and SMC_I3(OUT1, D1, S, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I8(shcheckCKD1lh, S, SE_bar);

    and SMC_I9(shcheckCKD2lh, S_bar, SE_bar);

    buf SMC_I10(shcheckCKSDlh, SE);

    not SMC_I11(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFMQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFMQM8RA (D1, D2, S, SD, SE, CK, Q);
  input D1, D2, S, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(S_bar, S);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT0, D2, S_bar, SE_bar);
    and SMC_I3(OUT1, D1, S, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I8(shcheckCKD1lh, S, SE_bar);

    and SMC_I9(shcheckCKD2lh, S_bar, SE_bar);

    buf SMC_I10(shcheckCKSDlh, SE);

    not SMC_I11(shcheckCKSlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D2 )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge S, posedge CK &&&
        (shcheckCKSlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D1, posedge CK &&&
        (shcheckCKD1lh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D2, posedge CK &&&
        (shcheckCKD2lh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), negedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), negedge D2, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), negedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSlh === 1'b1), posedge S, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD1lh === 1'b1), posedge D1, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKD2lh === 1'b1), posedge D2, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFMQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBM1RA (D, SD, SE, CK, QB);
  input D, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBM2RA (D, SD, SE, CK, QB);
  input D, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBM4RA (D, SD, SE, CK, QB);
  input D, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBM8RA (D, SD, SE, CK, QB);
  input D, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(shcheckCKDlh, SE);

    buf SMC_I5(shcheckCKSDlh, SE);


  specify


    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBRM1RA (D, RB, SD, SE, CK, QB);
  input D, RB, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBRM2RA (D, RB, SD, SE, CK, QB);
  input D, RB, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBRM4RA (D, RB, SD, SE, CK, QB);
  input D, RB, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQBRM8RA (D, RB, SD, SE, CK, QB);
  input D, RB, SD, SE, CK;
  output QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I4(SE_bar, SE);
    and SMC_I5(shcheckCKDlh, RB, SE_bar);

    and SMC_I6(shcheckCKSDlh, RB, SE);

    buf SMC_I7(shcheckCKSElh, RB);


  specify


    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQBRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQM1RA (D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(shcheckCKDlh, SE);

    buf SMC_I4(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);


    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQM2RA (D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(shcheckCKDlh, SE);

    buf SMC_I4(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);


    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQM4RA (D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(shcheckCKDlh, SE);

    buf SMC_I4(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);


    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQM8RA (D, SD, SE, CK, Q);
  input D, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(shcheckCKDlh, SE);

    buf SMC_I4(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);


    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRM1RA (D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, RB, SE_bar);

    and SMC_I5(shcheckCKSDlh, RB, SE);

    buf SMC_I6(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRM2RA (D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, RB, SE_bar);

    and SMC_I5(shcheckCKSDlh, RB, SE);

    buf SMC_I6(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRM4RA (D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, RB, SE_bar);

    and SMC_I5(shcheckCKSDlh, RB, SE);

    buf SMC_I6(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRM8RA (D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, RB, SE_bar);

    and SMC_I5(shcheckCKSDlh, RB, SE);

    buf SMC_I6(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRSM1RA (D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I5(shcheckCKRBlh, SB);

    buf SMC_I6(shcheckCKSBlh, RB);

    and SMC_I7(shcheckCKSDlh, RB, SB, SE);

    and SMC_I8(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRSM2RA (D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I5(shcheckCKRBlh, SB);

    buf SMC_I6(shcheckCKSBlh, RB);

    and SMC_I7(shcheckCKSDlh, RB, SB, SE);

    and SMC_I8(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRSM4RA (D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I5(shcheckCKRBlh, SB);

    buf SMC_I6(shcheckCKSBlh, RB);

    and SMC_I7(shcheckCKSDlh, RB, SB, SE);

    and SMC_I8(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQRSM8RA (D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I5(shcheckCKRBlh, SB);

    buf SMC_I6(shcheckCKSBlh, RB);

    and SMC_I7(shcheckCKSDlh, RB, SB, SE);

    and SMC_I8(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQSM1RA (D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, SB, SE_bar);

    and SMC_I5(shcheckCKSDlh, SB, SE);

    buf SMC_I6(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQSM2RA (D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, SB, SE_bar);

    and SMC_I5(shcheckCKSDlh, SB, SE);

    buf SMC_I6(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQSM4RA (D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, SB, SE_bar);

    and SMC_I5(shcheckCKSDlh, SB, SE);

    buf SMC_I6(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQSM8RA (D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    mux21 SMC_I0(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I1(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I2(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I3(SE_bar, SE);
    and SMC_I4(shcheckCKDlh, SB, SE_bar);

    and SMC_I5(shcheckCKSDlh, SB, SE);

    buf SMC_I6(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZRM1RA (D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, D, RB, SE_bar);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    not SMC_I7(shcheckCKRBlh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZRM2RA (D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, D, RB, SE_bar);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    not SMC_I7(shcheckCKRBlh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZRM4RA (D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, D, RB, SE_bar);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    not SMC_I7(shcheckCKRBlh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZRM8RA (D, RB, SD, SE, CK, Q);
  input D, RB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, D, RB, SE_bar);
    or SMC_I3(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I4(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I5(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I6(shcheckCKDlh, SE);

    not SMC_I7(shcheckCKRBlh, SE);

    buf SMC_I8(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZRSM1RA (D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SB_bar, SB);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT0, RB, SB_bar, SE_bar);
    and SMC_I3(OUT1, D, RB, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I8(shcheckCKDlh, RB, SE_bar);

    not SMC_I9(shcheckCKRBlh, SE);

    and SMC_I10(shcheckCKSBlh, RB, SE_bar);

    buf SMC_I11(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZRSM2RA (D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SB_bar, SB);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT0, RB, SB_bar, SE_bar);
    and SMC_I3(OUT1, D, RB, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I8(shcheckCKDlh, RB, SE_bar);

    not SMC_I9(shcheckCKRBlh, SE);

    and SMC_I10(shcheckCKSBlh, RB, SE_bar);

    buf SMC_I11(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZRSM4RA (D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SB_bar, SB);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT0, RB, SB_bar, SE_bar);
    and SMC_I3(OUT1, D, RB, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I8(shcheckCKDlh, RB, SE_bar);

    not SMC_I9(shcheckCKRBlh, SE);

    and SMC_I10(shcheckCKSBlh, RB, SE_bar);

    buf SMC_I11(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZRSM8RA (D, RB, SB, SD, SE, CK, Q);
  input D, RB, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    not SMC_I0(SB_bar, SB);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT0, RB, SB_bar, SE_bar);
    and SMC_I3(OUT1, D, RB, SE_bar);
    and SMC_I4(OUT2, SD, SE);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I8(shcheckCKDlh, RB, SE_bar);

    not SMC_I9(shcheckCKRBlh, SE);

    and SMC_I10(shcheckCKSBlh, RB, SE_bar);

    buf SMC_I11(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZSM1RA (D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, D, SE_bar);
    not SMC_I3(SB_bar, SB);
    and SMC_I4(OUT2, SB_bar, SE_bar);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(shcheckCKDlh, SE);

    not SMC_I9(shcheckCKSBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZSM2RA (D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, D, SE_bar);
    not SMC_I3(SB_bar, SB);
    and SMC_I4(OUT2, SB_bar, SE_bar);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(shcheckCKDlh, SE);

    not SMC_I9(shcheckCKSBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZSM4RA (D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, D, SE_bar);
    not SMC_I3(SB_bar, SB);
    and SMC_I4(OUT2, SB_bar, SE_bar);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(shcheckCKDlh, SE);

    not SMC_I9(shcheckCKSBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFQZSM8RA (D, SB, SD, SE, CK, Q);
  input D, SB, SD, SE, CK;
  output Q;
  reg notifier;

  wire SMC_NS_IN;
    and SMC_I0(OUT0, SD, SE);
    not SMC_I1(SE_bar, SE);
    and SMC_I2(OUT1, D, SE_bar);
    not SMC_I3(SB_bar, SB);
    and SMC_I4(OUT2, SB_bar, SE_bar);
    or SMC_I5(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I6(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I7(Q, SMC_IQ);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(shcheckCKDlh, SE);

    not SMC_I9(shcheckCKSBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFQZSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRM1RA (D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SE_bar);

    and SMC_I7(shcheckCKSDlh, RB, SE);

    buf SMC_I8(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRM2RA (D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SE_bar);

    and SMC_I7(shcheckCKSDlh, RB, SE);

    buf SMC_I8(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRM4RA (D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SE_bar);

    and SMC_I7(shcheckCKSDlh, RB, SE);

    buf SMC_I8(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRM8RA (D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SE_bar);

    and SMC_I7(shcheckCKSDlh, RB, SE);

    buf SMC_I8(shcheckCKSElh, RB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge RB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge RB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (RB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (RB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (RB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (RB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (RB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (RB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (RB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (RB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (RB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery RB-lh CK-lh ()
    $recovery(posedge RB, posedge CK, 0.0, notifier);

    // removal RB-lh CK-lh ()
    $hold(posedge CK, posedge RB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw RB-hl NS-hl ()
    $width(negedge RB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRSM1RA (D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I7(shcheckCKRBlh, SB);

    buf SMC_I8(shcheckCKSBlh, RB);

    and SMC_I9(shcheckCKSDlh, RB, SB, SE);

    and SMC_I10(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRSM2RA (D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I7(shcheckCKRBlh, SB);

    buf SMC_I8(shcheckCKSBlh, RB);

    and SMC_I9(shcheckCKSDlh, RB, SB, SE);

    and SMC_I10(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRSM4RA (D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I7(shcheckCKRBlh, SB);

    buf SMC_I8(shcheckCKSBlh, RB);

    and SMC_I9(shcheckCKSDlh, RB, SB, SE);

    and SMC_I10(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFRSM8RA (D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;


    inv_clr0 SMC_I0(.qn(SMC_IQN), .clr(RB), .pre(SB), .inp(SMC_IQ)
          );
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB) );

  `else // functional //

    dff_p0 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(RB),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, RB, SB, SE_bar);

    buf SMC_I7(shcheckCKRBlh, SB);

    buf SMC_I8(shcheckCKSBlh, RB);

    and SMC_I9(shcheckCKSDlh, RB, SB, SE);

    and SMC_I10(shcheckCKSElh, RB, SB);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc RB --> Q
    (negedge RB => ( Q +: D )) = (0.0, 0.0);

    // arc RB --> QB
    (negedge RB => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK &&&
        (shcheckCKSElh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSElh === 1'b1), posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge RB, 0.0, notifier );

    // recovery
    $recovery( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // recovery
    $recovery( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // removal
    $hold( posedge RB, posedge SB, 0.0, notifier );

    // removal
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // removal
    $hold( posedge SB, posedge RB, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge RB, 0.0, 0, notifier );

    // mpw
    $width( negedge SB, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFSM1RA (D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, SB, SE_bar);

    and SMC_I7(shcheckCKSDlh, SB, SE);

    buf SMC_I8(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFSM2RA (D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, SB, SE_bar);

    and SMC_I7(shcheckCKSDlh, SB, SE);

    buf SMC_I8(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFSM4RA (D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, SB, SE_bar);

    and SMC_I7(shcheckCKSDlh, SB, SE);

    buf SMC_I8(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFSM8RA (D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    mux21 SMC_I1(SMC_NS_IN, SD, D, SE);

  `ifdef functional // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB) );

  `else // functional //

    dff_p1 SMC_I2(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(SB), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I3(Q, SMC_IQ);

    buf SMC_I4(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I5(SE_bar, SE);
    and SMC_I6(shcheckCKDlh, SB, SE_bar);

    and SMC_I7(shcheckCKSDlh, SB, SE);

    buf SMC_I8(shcheckCKSElh, SB);


  specify


    // arc CK --> Q
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);

    // arc SB --> Q
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( Q +: D )) = (0.0, 0.0);

    // arc SB --> QB
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b0 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b0 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b0 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b0)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    if (CK===1'b1 && D===1'b1 && SD===1'b1 && SE===1'b1)
        (negedge SB => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (negedge SB => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (SB&!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (SB&!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh (SB)
    $setup(negedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SE-lh CK-lh (SB)
    $setup(posedge SE &&& (shcheckCKSElh === 1'b1),
        posedge CK &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // setup SD-hl CK-lh (SB&SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SB&SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (SB&!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        negedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SE-lh CK-lh (SB)
    $hold(posedge CK &&& (shcheckCKSElh === 1'b1),
        posedge SE &&& (shcheckCKSElh === 1'b1), 0.0, notifier);

    // hold SD-hl CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SB&SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // recovery SB-lh CK-lh ()
    $recovery(posedge SB, posedge CK, 0.0, notifier);

    // removal SB-lh CK-lh ()
    $hold(posedge CK, posedge SB, 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    // mpw SB-hl NS-hl ()
    $width(negedge SB, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRM1RA (D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, RB, SE_bar);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(shcheckCKDlh, SE);

    not SMC_I9(shcheckCKRBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
       (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRM2RA (D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, RB, SE_bar);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(shcheckCKDlh, SE);

    not SMC_I9(shcheckCKRBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
       (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRM4RA (D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, RB, SE_bar);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(shcheckCKDlh, SE);

    not SMC_I9(shcheckCKRBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
       (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRM8RA (D, RB, SD, SE, CK, Q, QB);
  input D, RB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, RB, SE_bar);
    or SMC_I4(SMC_NS_IN, OUT0, OUT1);


  `ifdef functional // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I5(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I6(Q, SMC_IQ);

    buf SMC_I7(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I8(shcheckCKDlh, SE);

    not SMC_I9(shcheckCKRBlh, SE);

    buf SMC_I10(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
       (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( Q +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b0 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b0 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b1 && SE===1'b1)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b1 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b0 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    if (D===1'b1 && RB===1'b1 && SD===1'b0 && SE===1'b0)
        (posedge CK => ( QB +: D )) = (0.0, 0.0);
    ifnone
        (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup D-hl CK-lh (!SE)
    $setup(negedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup D-lh CK-lh (!SE)
    $setup(posedge D &&& (shcheckCKDlh === 1'b1),
        posedge CK &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // setup RB-hl CK-lh (!SE)
    $setup(negedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup RB-lh CK-lh (!SE)
    $setup(posedge RB &&& (shcheckCKRBlh === 1'b1),
        posedge CK &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // setup SE-hl CK-lh ()
    $setup(negedge SE, posedge CK, 0.0, notifier);

    // setup SE-lh CK-lh ()
    $setup(posedge SE, posedge CK, 0.0, notifier);

    // setup SD-hl CK-lh (SE)
    $setup(negedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // setup SD-lh CK-lh (SE)
    $setup(posedge SD &&& (shcheckCKSDlh === 1'b1),
        posedge CK &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold D-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        negedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold D-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKDlh === 1'b1),
        posedge D &&& (shcheckCKDlh === 1'b1), 0.0, notifier);

    // hold RB-hl CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        negedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold RB-lh CK-lh (!SE)
    $hold(posedge CK &&& (shcheckCKRBlh === 1'b1),
        posedge RB &&& (shcheckCKRBlh === 1'b1), 0.0, notifier);

    // hold SE-hl CK-lh ()
    $hold(posedge CK, negedge SE, 0.0, notifier);

    // hold SE-lh CK-lh ()
    $hold(posedge CK, posedge SE, 0.0, notifier);

    // hold SD-hl CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        negedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // hold SD-lh CK-lh (SE)
    $hold(posedge CK &&& (shcheckCKSDlh === 1'b1),
        posedge SD &&& (shcheckCKSDlh === 1'b1), 0.0, notifier);

    // mpw CK-lh NS-lh ()
    $width(posedge CK, 0.0, 0, notifier);

    // mpw CK-hl NS-hl ()
    $width(negedge CK, 0.0, 0, notifier);

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRSM1RA (D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(SB_bar, SB);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT0, RB, SB_bar, SE_bar);
    and SMC_I4(OUT1, D, RB, SE_bar);
    and SMC_I5(OUT2, SD, SE);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I10(shcheckCKDlh, RB, SE_bar);

    not SMC_I11(shcheckCKRBlh, SE);

    and SMC_I12(shcheckCKSBlh, RB, SE_bar);

    buf SMC_I13(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRSM2RA (D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(SB_bar, SB);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT0, RB, SB_bar, SE_bar);
    and SMC_I4(OUT1, D, RB, SE_bar);
    and SMC_I5(OUT2, SD, SE);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I10(shcheckCKDlh, RB, SE_bar);

    not SMC_I11(shcheckCKRBlh, SE);

    and SMC_I12(shcheckCKSBlh, RB, SE_bar);

    buf SMC_I13(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRSM4RA (D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(SB_bar, SB);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT0, RB, SB_bar, SE_bar);
    and SMC_I4(OUT1, D, RB, SE_bar);
    and SMC_I5(OUT2, SD, SE);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I10(shcheckCKDlh, RB, SE_bar);

    not SMC_I11(shcheckCKRBlh, SE);

    and SMC_I12(shcheckCKSBlh, RB, SE_bar);

    buf SMC_I13(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZRSM8RA (D, RB, SB, SD, SE, CK, Q, QB);
  input D, RB, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    not SMC_I1(SB_bar, SB);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT0, RB, SB_bar, SE_bar);
    and SMC_I4(OUT1, D, RB, SE_bar);
    and SMC_I5(OUT2, SD, SE);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    and SMC_I10(shcheckCKDlh, RB, SE_bar);

    not SMC_I11(shcheckCKRBlh, SE);

    and SMC_I12(shcheckCKSBlh, RB, SE_bar);

    buf SMC_I13(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( negedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge RB, posedge CK &&&
        (shcheckCKRBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), negedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKRBlh === 1'b1), posedge RB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZRSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZSM1RA (D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, SE_bar);
    not SMC_I4(SB_bar, SB);
    and SMC_I5(OUT2, SB_bar, SE_bar);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I10(shcheckCKDlh, SE);

    not SMC_I11(shcheckCKSBlh, SE);

    buf SMC_I12(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZSM1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZSM2RA (D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, SE_bar);
    not SMC_I4(SB_bar, SB);
    and SMC_I5(OUT2, SB_bar, SE_bar);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I10(shcheckCKDlh, SE);

    not SMC_I11(shcheckCKSBlh, SE);

    buf SMC_I12(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZSM2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZSM4RA (D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, SE_bar);
    not SMC_I4(SB_bar, SB);
    and SMC_I5(OUT2, SB_bar, SE_bar);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I10(shcheckCKDlh, SE);

    not SMC_I11(shcheckCKSBlh, SE);

    buf SMC_I12(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZSM4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module SDFZSM8RA (D, SB, SD, SE, CK, Q, QB);
  input D, SB, SD, SE, CK;
  output Q, QB;
  reg notifier;

    not SMC_I0(SMC_IQN, SMC_IQ);
  wire SMC_NS_IN;
    and SMC_I1(OUT0, SD, SE);
    not SMC_I2(SE_bar, SE);
    and SMC_I3(OUT1, D, SE_bar);
    not SMC_I4(SB_bar, SB);
    and SMC_I5(OUT2, SB_bar, SE_bar);
    or SMC_I6(SMC_NS_IN, OUT0, OUT1, OUT2);


  `ifdef functional // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1) );

  `else // functional //

    dff_p0 SMC_I7(.q(SMC_IQ), .d(SMC_NS_IN), .clk(CK), .clear(1'b1),
          .preset(1'b1), .notifier(notifier) );

  `endif // functional //

    //  output pins

    buf SMC_I8(Q, SMC_IQ);

    buf SMC_I9(QB, SMC_IQN);


  `ifdef functional // functional //

  `else // functional //
    not SMC_I10(shcheckCKDlh, SE);

    not SMC_I11(shcheckCKSBlh, SE);

    buf SMC_I12(shcheckCKSDlh, SE);


  specify


    // arc CK --> Q
    (posedge CK => ( Q +: D )) = (0.0, 0.0);

    // arc CK --> QB
    (posedge CK => ( QB +: D )) = (0.0, 0.0);



    // setup
    $setup( posedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge D, posedge CK &&&
        (shcheckCKDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SD, posedge CK &&&
        (shcheckCKSDlh === 1'b1), 0.0, notifier );

    // setup
    $setup( posedge SE, posedge CK, 0.0, notifier );

    // setup
    $setup( posedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // setup
    $setup( negedge SB, posedge CK &&&
        (shcheckCKSBlh === 1'b1), 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), posedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), negedge D, 0.0, notifier );

    // hold
    $hold( posedge CK, negedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKDlh === 1'b1), posedge D, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSDlh === 1'b1), negedge SD, 0.0, notifier );

    // hold
    $hold( posedge CK, posedge SE, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), posedge SB, 0.0, notifier );

    // hold
    $hold( posedge CK &&&
        (shcheckCKSBlh === 1'b1), negedge SB, 0.0, notifier );

    // mpw
    $width( negedge CK, 0.0, 0, notifier );

    // mpw
    $width( posedge CK, 0.0, 0, notifier );

    $period( posedge CK, 0, notifier );
    $period( negedge CK, 0, notifier );

  endspecify

  `endif // functional //
endmodule     // SDFZSM8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module TIE0R (Z);
  output Z;

    buf SMC_I0(Z, 1'b0);


  `ifdef functional // functional //

  `else // functional //

  specify




  endspecify

  `endif // functional //
endmodule     // TIE0R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module TIE1R (Z);
  output Z;

    buf SMC_I0(Z, 1'b1);


  `ifdef functional // functional //

  `else // functional //

  specify




  endspecify

  `endif // functional //
endmodule     // TIE1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR2M0RA (A, B, Z);
  input A, B;
  output Z;

    xnor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR2M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR2M1RA (A, B, Z);
  input A, B;
  output Z;

    xnor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR2M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR2M2RA (A, B, Z);
  input A, B;
  output Z;

    xnor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR2M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR2M4RA (A, B, Z);
  input A, B;
  output Z;

    xnor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR2M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR2M6RA (A, B, Z);
  input A, B;
  output Z;

    xnor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR2M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR2M8RA (A, B, Z);
  input A, B;
  output Z;

    xnor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR2M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR3M0RA ( Z, A, B, C );
   input A, B, C;
   output Z;

    xnor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR3M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR3M1R ( Z, A, B, C );
   input A, B, C;
   output Z;

    xnor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR3M1R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR3M2R ( Z, A, B, C );
   input A, B, C;
   output Z;

    xnor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR3M2R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR3M4R ( Z, A, B, C );
   input A, B, C;
   output Z;

    xnor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR3M4R //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR3M6RA ( Z, A, B, C );
   input A, B, C;
   output Z;

    xnor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR3M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR3M8RA ( Z, A, B, C );
   input A, B, C;
   output Z;

    xnor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR3M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR4M1RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      XNR4_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR4M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR4M2RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      XNR4_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR4M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR4M4RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      XNR4_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR4M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XNR4M8RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      XNR4_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XNR4M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M0RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M1RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M2RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M3RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M3RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M4RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M6RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR2M8RA (A, B, Z);
  input A, B;
  output Z;

    xor SMC_I0(Z, A, B);


  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR2M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR3M0RA ( Z, A, B, C );
   input A, B, C;
   output Z;

   xor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR3M0RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR3M1RA ( Z, A, B, C );
   input A, B, C;
   output Z;

   xor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR3M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR3M2RA ( Z, A, B, C );
   input A, B, C;
   output Z;

   xor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR3M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR3M4RA ( Z, A, B, C );
   input A, B, C;
   output Z;

   xor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR3M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR3M6RA ( Z, A, B, C );
   input A, B, C;
   output Z;

   xor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR3M6RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR3M8RA ( Z, A, B, C );
   input A, B, C;
   output Z;

   xor (Z, A, B, C);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR3M8RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR4M1RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      XOR4_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR4M1RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR4M2RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      XOR4_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR4M2RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR4M4RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      XOR4_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR4M4RA //
`endcelldefine
`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif

`celldefine
module XOR4M8RA ( Z, A, B, C, D );
   input A, B, C, D;
   output Z;
      XOR4_UDP4(Z, A, B, C, D);

  `ifdef functional // functional //

  `else // functional //

  specify


    // arc A --> Z
    if (B===1'b0 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b0 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b0 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b0)
        (A => Z) = (0.0, 0.0);
    if (B===1'b1 && C===1'b1 && D===1'b1)
        (A => Z) = (0.0, 0.0);
    ifnone
        (A => Z) = (0.0, 0.0);

    // arc B --> Z
    if (A===1'b0 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b0 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b0 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b0)
        (B => Z) = (0.0, 0.0);
    if (A===1'b1 && C===1'b1 && D===1'b1)
        (B => Z) = (0.0, 0.0);
    ifnone
        (B => Z) = (0.0, 0.0);

    // arc C --> Z
    if (A===1'b0 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b0)
        (C => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && D===1'b1)
        (C => Z) = (0.0, 0.0);
    ifnone
        (C => Z) = (0.0, 0.0);

    // arc D --> Z
    if (A===1'b0 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b0 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b0 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b0)
        (D => Z) = (0.0, 0.0);
    if (A===1'b1 && B===1'b1 && C===1'b1)
        (D => Z) = (0.0, 0.0);
    ifnone
        (D => Z) = (0.0, 0.0);



  endspecify

  `endif // functional //
endmodule     // XOR4M8RA //
`endcelldefine

///////////////////////////////////////////////////////////////////////////


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AO31_UDP4(Z, A1, A2, A3, B);
output Z;
input A1, A2, A3, B;
table
// A1  A2  A3  B : Z
    ?   ?   ?  1  : 1;
    1   1   1  ?  : 1;
    ?   ?   0  0  : 0;
    ?   0   ?  0  : 0;
    0   ?   ?  0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AO32_UDP5(Z, A1, A2, A3, B1, B2);
output Z;
input A1, A2, A3, B1, B2;
table
// A1  A2  A3  B1  B2 : Z
    ?   ?   ?   1   1  : 1;
    1   1   1   ?   ?  : 1;
    0   ?   ?   ?   0  : 0;
    ?   ?   0   0   ?  : 0;
    0   ?   ?   0   ?  : 0;
    ?   ?   0   ?   0  : 0;
    ?   0   ?   0   ?  : 0;
    ?   0   ?   ?   0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AO33_UDP6(Z, A1, A2, A3, B1, B2, B3);
output Z;
input A1, A2, A3, B1, B2, B3;
table
// A1  A2  A3  B1  B2  B3 : Z
    ?   ?   ?   1   1   1  : 1;
    1   1   1   ?   ?   ?  : 1;
    0   ?   ?   0   ?   ?  : 0;
    ?   ?   0   ?   ?   0  : 0;
    0   ?   ?   ?   ?   0  : 0;
    ?   0   ?   0   ?   ?  : 0;
    ?   ?   0   ?   0   ?  : 0;
    ?   0   ?   ?   0   ?  : 0;
    ?   0   ?   ?   ?   0  : 0;
    ?   ?   0   0   ?   ?  : 0;
    0   ?   ?   ?   0   ?  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AO221_UDP5(Z, A1, A2, B1, B2, C);
output Z;
input A1, A2, B1, B2, C;
table
// A1  A2  B1  B2  C : Z
    ?   ?   ?   ?  1  : 1;
    ?   ?   1   1  ?  : 1;
    1   1   ?   ?  ?  : 1;
    ?   0   ?   0  0  : 0;
    ?   0   0   ?  0  : 0;
    0   ?   0   ?  0  : 0;
    0   ?   ?   0  0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive AO222_UDP6(Z, A1, A2, B1, B2, C1, C2);
output Z;
input A1, A2, B1, B2, C1, C2;
table
// A1  A2  B1  B2  C1  C2 : Z
    ?   ?   1   1   ?   ?  : 1;
    ?   ?   ?   ?   1   1  : 1;
    1   1   ?   ?   ?   ?  : 1;
    ?   0   ?   0   0   ?  : 0;
    0   ?   0   ?   ?   0  : 0;
    0   ?   0   ?   0   ?  : 0;
    ?   0   0   ?   0   ?  : 0;
    0   ?   ?   0   ?   0  : 0;
    0   ?   ?   0   0   ?  : 0;
    ?   0   0   ?   ?   0  : 0;
    ?   0   ?   0   ?   0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive DFEQZR_UDP__OUT__(__OUT__, D, E, IQ, RB);
output __OUT__;
input D, E, IQ, RB;
table
// D  E  IQ  RB : __OUT__
   ?  0   1   1  : 1;
   1  1   ?   1  : 1;
   0  1   ?   ?  : 0;
   ?  0   0   ?  : 0;
   ?  ?   ?   0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive DFEZR_UDP__OUT__(__OUT__, D, E, IQ, RB);
output __OUT__;
input D, E, IQ, RB;
table
// D  E  IQ  RB : __OUT__
   ?  0   1   1  : 1;
   1  1   ?   1  : 1;
   0  1   ?   ?  : 0;
   ?  0   0   ?  : 0;
   ?  ?   ?   0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MAO222_UDP3(Z, A, B, C);
output Z;
input A, B, C;
table
// A  B  C : Z
   1  ?  1  : 1;
   1  1  ?  : 1;
   ?  1  1  : 1;
   0  0  ?  : 0;
   0  ?  0  : 0;
   ?  0  0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MAOI2223_UDP4(Z, A, B, C, D);
output Z;
input A, B, C, D;
table
// A  B  C  D : Z
   ?  ?  0  0  : 1;
   ?  0  ?  0  : 1;
   0  0  0  ?  : 1;
   0  ?  ?  0  : 1;
   ?  ?  1  1  : 0;
   1  ?  ?  1  : 0;
   1  1  1  ?  : 0;
   ?  1  ?  1  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MAOI222_UDP3(Z, A, B, C);
output Z;
input A, B, C;
table
// A  B  C : Z
   0  0  ?  : 1;
   0  ?  0  : 1;
   ?  0  0  : 1;
   1  ?  1  : 0;
   1  1  ?  : 0;
   ?  1  1  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MOAI22_UDP4(Z, A1, A2, B1, B2);
output Z;
input A1, A2, B1, B2;
table
// A1  A2  B1  B2 : Z
    ?   ?   1   1  : 1;
    0   0   ?   ?  : 1;
    ?   1   0   ?  : 0;
    1   ?   ?   0  : 0;
    1   ?   0   ?  : 0;
    ?   1   ?   0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OA211_UDP4(Z, A1, A2, B, C);
output Z;
input A1, A2, B, C;
table
// A1  A2  B  C : Z
    ?   1  1  1  : 1;
    1   ?  1  1  : 1;
    ?   ?  ?  0  : 0;
    0   0  ?  ?  : 0;
    ?   ?  0  ?  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OA221_UDP5(Z, A1, A2, B1, B2, C);
output Z;
input A1, A2, B1, B2, C;
table
// A1  A2  B1  B2  C : Z
    ?   1   1   ?  1  : 1;
    ?   1   ?   1  1  : 1;
    1   ?   ?   1  1  : 1;
    1   ?   1   ?  1  : 1;
    ?   ?   ?   ?  0  : 0;
    ?   ?   0   0  ?  : 0;
    0   0   ?   ?  ?  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive OA222_UDP6(Z, A1, A2, B1, B2, C1, C2);
output Z;
input A1, A2, B1, B2, C1, C2;
table
// A1  A2  B1  B2  C1  C2 : Z
    1   ?   1   ?   1   ?  : 1;
    1   ?   ?   1   ?   1  : 1;
    ?   1   1   ?   ?   1  : 1;
    1   ?   ?   1   1   ?  : 1;
    1   ?   1   ?   ?   1  : 1;
    ?   1   ?   1   1   ?  : 1;
    ?   1   ?   1   ?   1  : 1;
    ?   1   1   ?   1   ?  : 1;
    ?   ?   ?   ?   0   0  : 0;
    0   0   ?   ?   ?   ?  : 0;
    ?   ?   0   0   ?   ?  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive SDFE_UDP__OUT__(__OUT__, D, E, IQ, SD, SE);
output __OUT__;
input D, E, IQ, SD, SE;
table
// D  E  IQ  SD  SE : __OUT__
   ?  ?   ?   1   1  : 1;
   ?  0   1   ?   0  : 1;
   1  1   ?   ?   0  : 1;
   0  1   ?   ?   0  : 0;
   ?  ?   ?   0   1  : 0;
   ?  0   0   ?   0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive SDFEQB_UDP__OUT__(__OUT__, D, E, IQ, SD, SE);
output __OUT__;
input D, E, IQ, SD, SE;
table
// D  E  IQ  SD  SE : __OUT__
   ?  ?   ?   1   1  : 1;
   ?  0   1   ?   0  : 1;
   1  1   ?   ?   0  : 1;
   0  1   ?   ?   0  : 0;
   ?  ?   ?   0   1  : 0;
   ?  0   0   ?   0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive SDFEQ_UDP__OUT__(__OUT__, D, E, IQ, SD, SE);
output __OUT__;
input D, E, IQ, SD, SE;
table
// D  E  IQ  SD  SE : __OUT__
   ?  ?   ?   1   1  : 1;
   ?  0   1   ?   0  : 1;
   1  1   ?   ?   0  : 1;
   0  1   ?   ?   0  : 0;
   ?  ?   ?   0   1  : 0;
   ?  0   0   ?   0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive SDFEQR_UDP__OUT__(__OUT__, D, E, IQ, SD, SE);
output __OUT__;
input D, E, IQ, SD, SE;
table
// D  E  IQ  SD  SE : __OUT__
   ?  ?   ?   1   1  : 1;
   ?  0   1   ?   0  : 1;
   1  1   ?   ?   0  : 1;
   0  1   ?   ?   0  : 0;
   ?  ?   ?   0   1  : 0;
   ?  0   0   ?   0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive SDFEQZR_UDP__OUT__(__OUT__, D, E, IQ, RB, SD, SE);
output __OUT__;
input D, E, IQ, RB, SD, SE;
table
// D  E  IQ  RB  SD  SE : __OUT__
   1  1   ?   1   ?   0  : 1;
   ?  ?   ?   ?   1   1  : 1;
   ?  0   1   1   ?   0  : 1;
   ?  ?   ?   0   ?   0  : 0;
   ?  0   0   ?   ?   0  : 0;
   0  1   ?   ?   ?   0  : 0;
   ?  ?   ?   ?   0   1  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive SDFER_UDP__OUT__(__OUT__, D, E, IQ, SD, SE);
output __OUT__;
input D, E, IQ, SD, SE;
table
// D  E  IQ  SD  SE : __OUT__
   ?  ?   ?   1   1  : 1;
   ?  0   1   ?   0  : 1;
   1  1   ?   ?   0  : 1;
   0  1   ?   ?   0  : 0;
   ?  ?   ?   0   1  : 0;
   ?  0   0   ?   0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive SDFEZR_UDP__OUT__(__OUT__, D, E, IQ, RB, SD, SE);
output __OUT__;
input D, E, IQ, RB, SD, SE;
table
// D  E  IQ  RB  SD  SE : __OUT__
   1  1   ?   1   ?   0  : 1;
   ?  ?   ?   ?   1   1  : 1;
   ?  0   1   1   ?   0  : 1;
   ?  ?   ?   0   ?   0  : 0;
   ?  0   0   ?   ?   0  : 0;
   0  1   ?   ?   ?   0  : 0;
   ?  ?   ?   ?   0   1  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive XNR4_UDP4(Z, A, B, C, D);
output Z;
input A, B, C, D;
table
// A  B  C  D : Z
   0  0  1  1  : 1;
   0  0  0  0  : 1;
   0  1  1  0  : 1;
   1  1  1  1  : 1;
   1  0  1  0  : 1;
   1  0  0  1  : 1;
   0  1  0  1  : 1;
   1  1  0  0  : 1;
   0  1  1  1  : 0;
   1  0  0  0  : 0;
   0  0  0  1  : 0;
   1  1  0  1  : 0;
   1  1  1  0  : 0;
   1  0  1  1  : 0;
   0  0  1  0  : 0;
   0  1  0  0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive XOR4_UDP4(Z, A, B, C, D);
output Z;
input A, B, C, D;
table
// A  B  C  D : Z
   0  1  1  1  : 1;
   1  0  0  0  : 1;
   0  0  0  1  : 1;
   1  1  0  1  : 1;
   1  1  1  0  : 1;
   1  0  1  1  : 1;
   0  0  1  0  : 1;
   0  1  0  0  : 1;
   0  0  1  1  : 0;
   0  0  0  0  : 0;
   0  1  1  0  : 0;
   1  1  1  1  : 0;
   1  0  1  0  : 0;
   1  0  0  1  : 0;
   0  1  0  1  : 0;
   1  1  0  0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive BEMXB_UDP5(PB, M0, M1, OA1, OA2, Z);
output PB;
input M0, M1, OA1, OA2, Z;
table
// M0  M1  OA1  OA2  Z : PB
    ?   1    1    ?  0  : 1;
    1   ?    1    ?  1  : 1;
    0   ?    ?    1  1  : 1;
    ?   0    ?    1  0  : 1;
    ?   1    0    ?  0  : 0;
    ?   0    ?    0  0  : 0;
    1   ?    0    ?  1  : 0;
    0   ?    ?    0  1  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive BEMX_UDP5(P, M0, M1, OA1, OA2, Z);
output P;
input M0, M1, OA1, OA2, Z;
table
// M0  M1  OA1  OA2  Z : P
    ?   1    0    ?  0  : 1;
    ?   0    ?    0  0  : 1;
    1   ?    0    ?  1  : 1;
    0   ?    ?    0  1  : 1;
    ?   1    1    ?  0  : 0;
    1   ?    1    ?  1  : 0;
    0   ?    ?    1  1  : 0;
    ?   0    ?    1  0  : 0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MUX3_UDP5(Z, A, B, C, S0, S1);
output Z;
input A, B, C, S0, S1;
table
// A  B  C  S0  S1 : Z
   0  ?  ?  0  0  :  0;
   1  ?  ?  0  0  :  1;
   ?  0  ?  1  0  :  0;
   ?  1  ?  1  0  :  1;
   ?  ?  0  0  1  :  0;
   ?  ?  1  0  1  :  1;
   ?  ?  0  1  1  :  0;
   ?  ?  1  1  1  :  1;
   0  0  ?  x  0  :  0;
   1  1  ?  x  0  :  1;
   ?  ?  0  x  1  :  0;
   ?  ?  1  x  1  :  1;
   0  ?  0  0  x  :  0;
   1  ?  1  0  x  :  1;
   ?  0  0  1  x  :  0;
   ?  1  1  1  x  :  1;
   1  1  1  x  x  :  1;
   0  0  0  x  x  :  0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MUX4_UDP6(Z, A, B, C, D, S0, S1);
output Z;
input A, B, C, D, S0, S1;
table
// A  B  C  D  S0  S1 : Z
   0  ?  ?  ?  0  0  :  0;
   1  ?  ?  ?  0  0  :  1;
   ?  0  ?  ?  1  0  :  0;
   ?  1  ?  ?  1  0  :  1;
   ?  ?  0  ?  0  1  :  0;
   ?  ?  1  ?  0  1  :  1;
   ?  ?  ?  0  1  1  :  0;
   ?  ?  ?  1  1  1  :  1;
   0  0  ?  ?  x  0  :  0;
   1  1  ?  ?  x  0  :  1;
   ?  ?  0  0  x  1  :  0;
   ?  ?  1  1  x  1  :  1;
   0  ?  0  ?  0  x  :  0;
   1  ?  1  ?  0  x  :  1;
   ?  0  ?  0  1  x  :  0;
   ?  1  ?  1  1  x  :  1;
   1  1  1  1  x  x  :  1;
   0  0  0  0  x  x  :  0;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MXB3_UDP5(Z, A, B, C, S0, S1);
output Z;
input A, B, C, S0, S1;
table
// A  B  C  S0  S1 : Z
   0  ?  ?  0  0  :  1;
   1  ?  ?  0  0  :  0;
   ?  0  ?  1  0  :  1;
   ?  1  ?  1  0  :  0;
   ?  ?  0  0  1  :  1;
   ?  ?  1  0  1  :  0;
   ?  ?  0  1  1  :  1;
   ?  ?  1  1  1  :  0;
   0  0  ?  x  0  :  1;
   1  1  ?  x  0  :  0;
   ?  ?  0  x  1  :  1;
   ?  ?  1  x  1  :  0;
   0  ?  0  0  x  :  1;
   1  ?  1  0  x  :  0;
   ?  0  0  1  x  :  1;
   ?  1  1  1  x  :  0;
   1  1  1  x  x  :  0;
   0  0  0  x  x  :  1;

endtable
endprimitive


`timescale 1 ns / 1 ps

`ifdef functional
				// none
`else
	`define SMC_NFORCE 1 	// Flag to force output to x if notifer changes
`endif


primitive MXB4_UDP6(Z, A, B, C, D, S0, S1);
output Z;
input A, B, C, D, S0, S1;
table
// A  B  C  D  S0  S1 : Z
   0  ?  ?  ?  0  0  :  1;
   1  ?  ?  ?  0  0  :  0;
   ?  0  ?  ?  1  0  :  1;
   ?  1  ?  ?  1  0  :  0;
   ?  ?  0  ?  0  1  :  1;
   ?  ?  1  ?  0  1  :  0;
   ?  ?  ?  0  1  1  :  1;
   ?  ?  ?  1  1  1  :  0;
   0  0  ?  ?  x  0  :  1;
   1  1  ?  ?  x  0  :  0;
   ?  ?  0  0  x  1  :  1;
   ?  ?  1  1  x  1  :  0;
   0  ?  0  ?  0  x  :  1;
   1  ?  1  ?  0  x  :  0;
   ?  0  ?  0  1  x  :  1;
   ?  1  ?  1  1  x  :  0;
   1  1  1  1  x  x  :  0;
   0  0  0  0  x  x  :  1;

endtable
endprimitive

// CR default primitives
// All cells assume preset and clear are active low


///////////////////////////////////////////////////////////////////////////
// This dff cell has a reset priority over preset

primitive udp_dff_p0(q, d, clk, clear, preset, notifier);
	output q;
	input  clk, clear, d, preset, notifier;
	reg q; /* declaring output as reg*/

	table
	// d  clk  clear  preset  notifier : state : q
           0   r    ?      1     ?    : ?  :  0  ; // clock in 0
           1   r    1      ?     ?    : ?  :  1  ; // clock in 1

           1   *    1      ?     ?    : 1  :  1  ; // reduce pessimism
           0   *    ?      1     ?    : 0  :  0  ; // reduce pessimism

           ?   f    ?      ?     ?    : ?  :  -  ; // no changes on negedge clk
           *   b    ?      ?     ?    : ?  :  -  ; // no changes when in switches

           ?   ?    0      ?     ?    : ?  :  0  ; // reset output; dominate

           ?   b    1      *     ?    : 1  :  1  ; // cover all transistions on set_
           1   x    1      *     ?    : 1  :  1  ; // cover all transistions on set_

           ?   ?    1      0     ?    : ?  :  1  ; // set output

           ?   b    *      1     ?    : 0  :  0  ; // cover all transistions on clr_
           0   x    *      1     ?    : 0  :  0  ; // cover all transistions on clr_

`ifdef SMC_NFORCE
	   ?   ?     ?      ?        *     :   ?   : x ;  // on any notifier event output x
`else
	   ?   ?     ?      ?        *     :   ?   : - ;  // ignore notifier changes in functional mode
`endif
	endtable
endprimitive

module dff_p0(q, d, clk, clear, preset, notifier);
   output q;
   input  clk, clear, d, preset, notifier;

   udp_dff_p0 D1(q, d, clk, clear, preset, notifier);
endmodule // dff_p0

///////////////////////////////////////////////////////////////////////////
// This cell has a preset priority over reset

primitive udp_dff_p1(q, d, clk, clear, preset, notifier);
	output q;
	input  clk, clear, d, preset, notifier;
	reg q; /* declaring output as reg*/

	table
	// d  clk  clear  preset  notifier : state : q
           0   r    ?      1     ?    : ?  :  0  ; // clock in 0
           1   r    1      ?     ?    : ?  :  1  ; // clock in 1

           1   *    1      ?     ?    : 1  :  1  ; // reduce pessimism
           0   *    ?      1     ?    : 0  :  0  ; // reduce pessimism

           ?   f    ?      ?     ?    : ?  :  -  ; // no changes on negedge clk
           *   b    ?      ?     ?    : ?  :  -  ; // no changes when in switches

           ?   ?    ?      0     ?    : ?  :  1  ; // set output; dominate

           ?   b    1      *     ?    : 1  :  1  ; // cover all transistions on set_
           1   x    1      *     ?    : 1  :  1  ; // cover all transistions on set_

           ?   ?    0      1     ?    : ?  :  0  ; // reset output

           ?   b    *      1     ?    : 0  :  0  ; // cover all transistions on clr_
           0   x    *      1     ?    : 0  :  0  ; // cover all transistions on clr_
`ifdef SMC_NFORCE
	   ?   ?     ?      ?        *     :   ?   : x ;  // on any notifier event output x
`else
	   ?   ?     ?      ?        *     :   ?   : - ;  // ignore notifier changes in functional mode
`endif
	endtable
endprimitive

module dff_p1(q, d, clk, clear, preset, notifier);
   output q;
   input  clk, clear, d, preset, notifier;

   udp_dff_p1 D1(q, d, clk, clear, preset, notifier);
endmodule // dff_p1



///////////////////////////////////////////////////////////////////////////
//

primitive udp_inv_clr0 (qn, clr, pre, inp);
	output qn;
	input  clr, pre, inp;

	table

	//  	clr 	pre 	inp	: qn
		0	0	?	: 0;
		1	?	0	: 1;
		1	?	1	: 0;
		?	1	0	: 1;
		?	1	1	: 0;
		x	x	1	: 0;
		x	x	0	: 1;
	endtable
endprimitive

module inv_clr0 (qn, clr, pre, inp);
   output qn;
   input  clr, pre, inp;

   udp_inv_clr0 (qn, clr, pre, inp);
endmodule // inv_clr0


///////////////////////////////////////////////////////////////////////////
//

primitive udp_mux21 (q, data1, data0, dselect);
    output q;
    input data1, data0, dselect;

// FUNCTION :  TWO TO ONE MULTIPLEXER
table
//data1 data0 dselect :   q
        0     0       ?   :   0 ;
        1     1       ?   :   1 ;

        0     ?       1   :   0 ;
        1     ?       1   :   1 ;

        ?     0       0   :   0 ;
        ?     1       0   :   1 ;
endtable
endprimitive


module mux21 (q, data1, data0, dselect);
   output q;
   input  data1, data0, dselect;

   udp_mux21 m1(q, data1, data0, dselect);
endmodule // mux21

///////////////////////////////////////////////////////////////////////////
//

primitive udp_ldlatch_p0(q, d, en, clear, preset, notifier);
	output q;
	input  d, en, clear, preset, notifier;
	reg q;

	table
	// d  en  clear	 preset	 notifier : state : q
           1  1    1     ?        ?       : ?  :  1  ; //
           0  1    ?     1        ?       : ?  :  0  ; //
           1  *    1     ?        ?       : 1  :  1  ; // reduce pessimism
           0  *    ?     1        ?       : 0  :  0  ; // reduce pessimism
           *  0    ?     ?        ?       : ?  :  -  ; // no changes when in switches

           ?  ?    0     ?        ?       : ?  :  0  ; // reset output : reset dominate

           ?  0    1     *        ?       : 1  :  1  ; // cover all transistions on set_
           1  ?    1     *        ?       : 1  :  1  ; // cover all transistions on set_

           ?  ?    1     0        ?       : ?  :  1  ; // set output

           ?  0    *     1        ?       : 0  :  0  ; // cover all transistions on clr_
           0  ?    *     1        ?       : 0  :  0  ; // cover all transistions on clr_
`ifdef SMC_NFORCE
	   ?  ?    ?     ?        *       : ?  :  x ;  // on any notifier event output x
`else
	   ?  ?    ?     ?        *       : ?  :  - ;  // ignore notifier changes in functional mode
`endif
	endtable
endprimitive

module ldlatch_p0(q, d, en, clear, preset, notifier);
   output q;
   input  clear, preset, d, en, notifier;

   udp_ldlatch_p0 P1 (q, d, en, clear, preset, notifier);
endmodule // ldlatch_p0

///////////////////////////////////////////////////////////////////////////
//

primitive udp_ldlatch_p1(q, d, en, clear, preset, notifier);
	output q;
	input  clear, preset, d, en, notifier;
	reg q;

	table
	// d  en  clear	 preset	 notifier : state : q
           1  1   1   ?   ?   : ?  :  1  ; //
           0  1   ?   1   ?   : ?  :  0  ; //
           1  *   1   ?   ?   : 1  :  1  ; // reduce pessimism
           0  *   ?   1   ?   : 0  :  0  ; // reduce pessimism
           *  0   ?   ?   ?   : ?  :  -  ; // no changes when in switches
           ?  ?   ?   0   ?   : ?  :  1  ; // set output
           ?  0   1   *   ?   : 1  :  1  ; // cover all transistions on set_
           1  ?   1   *   ?   : 1  :  1  ; // cover all transistions on set_
           ?  ?   0   1   ?   : ?  :  0  ; // reset output
           ?  0   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
           0  ?   *   1   ?   : 0  :  0  ; // cover all transistions on clr_
`ifdef SMC_NFORCE
	   ?   ?    ?      ?        *     :   ?   : x ;  // on any notifier event output x
`else
	   ?   ?    ?      ?        *     :   ?   : - ;  // ignore notifier changes in functional mode
`endif
	endtable
endprimitive

module ldlatch_p1(q, d, en, clear, preset, notifier);
   output q;
   input clear, preset, d, en, notifier;

   udp_ldlatch_p1 P1 (q, d, en, clear, preset, notifier);
endmodule // ldlatch_p1
