/**
    Add the code for your adc_analog module here

*/
