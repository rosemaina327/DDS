/**

    This module wraps the basic ADC and adds a test DAC
*/
